library ieee;use ieee.std_logic_1164.all;entity fir_cs isport (  clk, reset : in std_logic;  in_1_1 : in std_logic_vector(5 downto 0);  in_1_2 : in std_logic_vector(5 downto 0);  in_1_3 : in std_logic_vector(5 downto 0);  in_1_4 : in std_logic_vector(5 downto 0);  in_1_5 : in std_logic_vector(5 downto 0);  in_1_6 : in std_logic_vector(4 downto 0);  in_1_7 : in std_logic_vector(3 downto 0);  in_1_8 : in std_logic_vector(2 downto 0);  in_1_9 : in std_logic_vector(1 downto 0);  in_1_10 : in std_logic_vector(0 downto 0);  in_5_4 : in std_logic_vector(0 downto 0);  in_5_5 : in std_logic_vector(0 downto 0);  in_5_6 : in std_logic_vector(1 downto 0);  in_5_7 : in std_logic_vector(1 downto 0);  in_5_8 : in std_logic_vector(1 downto 0);  in_5_9 : in std_logic_vector(1 downto 0);  in_5_10 : in std_logic_vector(0 downto 0);  in_5_11 : in std_logic_vector(0 downto 0);  in_7_3 : in std_logic_vector(0 downto 0);  in_7_4 : in std_logic_vector(0 downto 0);  in_7_5 : in std_logic_vector(0 downto 0);  in_7_6 : in std_logic_vector(0 downto 0);  in_7_7 : in std_logic_vector(0 downto 0);  in_7_8 : in std_logic_vector(0 downto 0);  in_9_4 : in std_logic_vector(0 downto 0);  in_9_5 : in std_logic_vector(0 downto 0);  in_9_6 : in std_logic_vector(1 downto 0);  in_9_7 : in std_logic_vector(1 downto 0);  in_9_8 : in std_logic_vector(1 downto 0);  in_9_9 : in std_logic_vector(1 downto 0);  in_9_10 : in std_logic_vector(0 downto 0);  in_9_11 : in std_logic_vector(0 downto 0);  in_13_1 : in std_logic_vector(5 downto 0);  in_13_2 : in std_logic_vector(5 downto 0);  in_13_3 : in std_logic_vector(5 downto 0);  in_13_4 : in std_logic_vector(5 downto 0);  in_13_5 : in std_logic_vector(5 downto 0);  in_13_6 : in std_logic_vector(4 downto 0);  in_13_7 : in std_logic_vector(3 downto 0);  in_13_8 : in std_logic_vector(2 downto 0);  in_13_9 : in std_logic_vector(1 downto 0);  in_13_10 : in std_logic_vector(0 downto 0);  out_1 : out std_logic_vector(1 downto 0);  out_2 : out std_logic_vector(1 downto 0);  out_3 : out std_logic_vector(1 downto 0);  out_4 : out std_logic_vector(1 downto 0);  out_5 : out std_logic_vector(1 downto 0);  out_6 : out std_logic_vector(1 downto 0);  out_7 : out std_logic_vector(1 downto 0);  out_8 : out std_logic_vector(0 downto 0);  out_9 : out std_logic_vector(0 downto 0);  out_10 : out std_logic_vector(0 downto 0);  out_11 : out std_logic_vector(0 downto 0));end fir_cs;architecture generated of fir_cs iscomponent faport (in1, in2, in3 : in  std_logic;      outs, outc    : out std_logic);end component;component haport (in1, in2   : in  std_logic;      outs, outc : out std_logic);end component;component fa_nocport (in1, in2, in3 : in  std_logic;      outs          : out std_logic);end component;component ha_nocport (in1, in2 : in  std_logic;      outs     : out std_logic);end component;component dffport (clk, reset : in std_logic;      d : in  std_logic;      q : out std_logic);end component;signal cellin_1_1 : std_logic_vector(5 downto 0);signal cellin_1_2 : std_logic_vector(5 downto 0);signal cellin_1_3 : std_logic_vector(5 downto 0);signal cellin_1_4 : std_logic_vector(5 downto 0);signal cellin_1_5 : std_logic_vector(5 downto 0);signal cellin_1_6 : std_logic_vector(4 downto 0);signal cellin_1_7 : std_logic_vector(3 downto 0);signal cellin_1_8 : std_logic_vector(2 downto 0);signal cellin_1_9 : std_logic_vector(1 downto 0);signal cellin_1_10 : std_logic_vector(0 downto 0);signal cellin_2_1 : std_logic_vector(3 downto 0);signal cellin_2_2 : std_logic_vector(3 downto 0);signal cellin_2_3 : std_logic_vector(3 downto 0);signal cellin_2_4 : std_logic_vector(3 downto 0);signal cellin_2_5 : std_logic_vector(2 downto 0);signal cellin_2_6 : std_logic_vector(3 downto 0);signal cellin_2_7 : std_logic_vector(2 downto 0);signal cellin_2_8 : std_logic_vector(0 downto 0);signal cellin_2_9 : std_logic_vector(1 downto 0);signal cellin_2_10 : std_logic_vector(0 downto 0);signal cellin_3_1 : std_logic_vector(2 downto 0);signal cellin_3_2 : std_logic_vector(2 downto 0);signal cellin_3_3 : std_logic_vector(2 downto 0);signal cellin_3_4 : std_logic_vector(2 downto 0);signal cellin_3_5 : std_logic_vector(1 downto 0);signal cellin_3_6 : std_logic_vector(2 downto 0);signal cellin_3_7 : std_logic_vector(0 downto 0);signal cellin_3_8 : std_logic_vector(0 downto 0);signal cellin_3_9 : std_logic_vector(1 downto 0);signal cellin_3_10 : std_logic_vector(0 downto 0);signal cellin_4_1 : std_logic_vector(1 downto 0);signal cellin_4_2 : std_logic_vector(1 downto 0);signal cellin_4_3 : std_logic_vector(1 downto 0);signal cellin_4_4 : std_logic_vector(1 downto 0);signal cellin_4_5 : std_logic_vector(1 downto 0);signal cellin_4_6 : std_logic_vector(0 downto 0);signal cellin_4_7 : std_logic_vector(0 downto 0);signal cellin_4_8 : std_logic_vector(0 downto 0);signal cellin_4_9 : std_logic_vector(1 downto 0);signal cellin_4_10 : std_logic_vector(0 downto 0);signal cellin_5_1 : std_logic_vector(1 downto 0);signal cellin_5_2 : std_logic_vector(1 downto 0);signal cellin_5_3 : std_logic_vector(1 downto 0);signal cellin_5_4 : std_logic_vector(2 downto 0);signal cellin_5_5 : std_logic_vector(2 downto 0);signal cellin_5_6 : std_logic_vector(2 downto 0);signal cellin_5_7 : std_logic_vector(2 downto 0);signal cellin_5_8 : std_logic_vector(2 downto 0);signal cellin_5_9 : std_logic_vector(3 downto 0);signal cellin_5_10 : std_logic_vector(1 downto 0);signal cellin_5_11 : std_logic_vector(0 downto 0);signal cellin_6_1 : std_logic_vector(1 downto 0);signal cellin_6_2 : std_logic_vector(1 downto 0);signal cellin_6_3 : std_logic_vector(2 downto 0);signal cellin_6_4 : std_logic_vector(1 downto 0);signal cellin_6_5 : std_logic_vector(1 downto 0);signal cellin_6_6 : std_logic_vector(1 downto 0);signal cellin_6_7 : std_logic_vector(1 downto 0);signal cellin_6_8 : std_logic_vector(1 downto 0);signal cellin_6_9 : std_logic_vector(1 downto 0);signal cellin_6_10 : std_logic_vector(1 downto 0);signal cellin_6_11 : std_logic_vector(0 downto 0);signal cellin_7_1 : std_logic_vector(1 downto 0);signal cellin_7_2 : std_logic_vector(1 downto 0);signal cellin_7_3 : std_logic_vector(1 downto 0);signal cellin_7_4 : std_logic_vector(2 downto 0);signal cellin_7_5 : std_logic_vector(2 downto 0);signal cellin_7_6 : std_logic_vector(2 downto 0);signal cellin_7_7 : std_logic_vector(2 downto 0);signal cellin_7_8 : std_logic_vector(2 downto 0);signal cellin_7_9 : std_logic_vector(1 downto 0);signal cellin_7_10 : std_logic_vector(1 downto 0);signal cellin_7_11 : std_logic_vector(0 downto 0);signal cellin_8_1 : std_logic_vector(1 downto 0);signal cellin_8_2 : std_logic_vector(1 downto 0);signal cellin_8_3 : std_logic_vector(1 downto 0);signal cellin_8_4 : std_logic_vector(1 downto 0);signal cellin_8_5 : std_logic_vector(1 downto 0);signal cellin_8_6 : std_logic_vector(1 downto 0);signal cellin_8_7 : std_logic_vector(1 downto 0);signal cellin_8_8 : std_logic_vector(0 downto 0);signal cellin_8_9 : std_logic_vector(1 downto 0);signal cellin_8_10 : std_logic_vector(1 downto 0);signal cellin_8_11 : std_logic_vector(0 downto 0);signal cellin_9_1 : std_logic_vector(1 downto 0);signal cellin_9_2 : std_logic_vector(1 downto 0);signal cellin_9_3 : std_logic_vector(1 downto 0);signal cellin_9_4 : std_logic_vector(2 downto 0);signal cellin_9_5 : std_logic_vector(2 downto 0);signal cellin_9_6 : std_logic_vector(3 downto 0);signal cellin_9_7 : std_logic_vector(3 downto 0);signal cellin_9_8 : std_logic_vector(2 downto 0);signal cellin_9_9 : std_logic_vector(3 downto 0);signal cellin_9_10 : std_logic_vector(2 downto 0);signal cellin_9_11 : std_logic_vector(1 downto 0);signal cellin_10_1 : std_logic_vector(1 downto 0);signal cellin_10_2 : std_logic_vector(1 downto 0);signal cellin_10_3 : std_logic_vector(2 downto 0);signal cellin_10_4 : std_logic_vector(1 downto 0);signal cellin_10_5 : std_logic_vector(1 downto 0);signal cellin_10_6 : std_logic_vector(2 downto 0);signal cellin_10_7 : std_logic_vector(2 downto 0);signal cellin_10_8 : std_logic_vector(1 downto 0);signal cellin_10_9 : std_logic_vector(2 downto 0);signal cellin_10_10 : std_logic_vector(0 downto 0);signal cellin_10_11 : std_logic_vector(1 downto 0);signal cellin_11_1 : std_logic_vector(1 downto 0);signal cellin_11_2 : std_logic_vector(1 downto 0);signal cellin_11_3 : std_logic_vector(1 downto 0);signal cellin_11_4 : std_logic_vector(1 downto 0);signal cellin_11_5 : std_logic_vector(1 downto 0);signal cellin_11_6 : std_logic_vector(1 downto 0);signal cellin_11_7 : std_logic_vector(1 downto 0);signal cellin_11_8 : std_logic_vector(1 downto 0);signal cellin_11_9 : std_logic_vector(0 downto 0);signal cellin_11_10 : std_logic_vector(0 downto 0);signal cellin_11_11 : std_logic_vector(1 downto 0);signal cellin_12_1 : std_logic_vector(1 downto 0);signal cellin_12_2 : std_logic_vector(1 downto 0);signal cellin_12_3 : std_logic_vector(1 downto 0);signal cellin_12_4 : std_logic_vector(1 downto 0);signal cellin_12_5 : std_logic_vector(1 downto 0);signal cellin_12_6 : std_logic_vector(1 downto 0);signal cellin_12_7 : std_logic_vector(1 downto 0);signal cellin_12_8 : std_logic_vector(1 downto 0);signal cellin_12_9 : std_logic_vector(0 downto 0);signal cellin_12_10 : std_logic_vector(0 downto 0);signal cellin_12_11 : std_logic_vector(1 downto 0);signal cellin_13_1 : std_logic_vector(8 downto 0);signal cellin_13_2 : std_logic_vector(8 downto 0);signal cellin_13_3 : std_logic_vector(7 downto 0);signal cellin_13_4 : std_logic_vector(7 downto 0);signal cellin_13_5 : std_logic_vector(8 downto 0);signal cellin_13_6 : std_logic_vector(6 downto 0);signal cellin_13_7 : std_logic_vector(5 downto 0);signal cellin_13_8 : std_logic_vector(4 downto 0);signal cellin_13_9 : std_logic_vector(2 downto 0);signal cellin_13_10 : std_logic_vector(1 downto 0);signal cellin_13_11 : std_logic_vector(1 downto 0);signal cellin_14_1 : std_logic_vector(5 downto 0);signal cellin_14_2 : std_logic_vector(5 downto 0);signal cellin_14_3 : std_logic_vector(5 downto 0);signal cellin_14_4 : std_logic_vector(5 downto 0);signal cellin_14_5 : std_logic_vector(4 downto 0);signal cellin_14_6 : std_logic_vector(4 downto 0);signal cellin_14_7 : std_logic_vector(2 downto 0);signal cellin_14_8 : std_logic_vector(3 downto 0);signal cellin_14_9 : std_logic_vector(0 downto 0);signal cellin_14_10 : std_logic_vector(2 downto 0);signal cellin_14_11 : std_logic_vector(0 downto 0);signal cellin_15_1 : std_logic_vector(3 downto 0);signal cellin_15_2 : std_logic_vector(3 downto 0);signal cellin_15_3 : std_logic_vector(3 downto 0);signal cellin_15_4 : std_logic_vector(2 downto 0);signal cellin_15_5 : std_logic_vector(3 downto 0);signal cellin_15_6 : std_logic_vector(3 downto 0);signal cellin_15_7 : std_logic_vector(1 downto 0);signal cellin_15_8 : std_logic_vector(1 downto 0);signal cellin_15_9 : std_logic_vector(1 downto 0);signal cellin_15_10 : std_logic_vector(0 downto 0);signal cellin_15_11 : std_logic_vector(0 downto 0);signal cellin_16_1 : std_logic_vector(2 downto 0);signal cellin_16_2 : std_logic_vector(2 downto 0);signal cellin_16_3 : std_logic_vector(2 downto 0);signal cellin_16_4 : std_logic_vector(1 downto 0);signal cellin_16_5 : std_logic_vector(2 downto 0);signal cellin_16_6 : std_logic_vector(1 downto 0);signal cellin_16_7 : std_logic_vector(1 downto 0);signal cellin_16_8 : std_logic_vector(2 downto 0);signal cellin_16_9 : std_logic_vector(0 downto 0);signal cellin_16_10 : std_logic_vector(0 downto 0);signal cellin_16_11 : std_logic_vector(0 downto 0);signal cellin_17_1 : std_logic_vector(1 downto 0);signal cellin_17_2 : std_logic_vector(1 downto 0);signal cellin_17_3 : std_logic_vector(1 downto 0);signal cellin_17_4 : std_logic_vector(1 downto 0);signal cellin_17_5 : std_logic_vector(1 downto 0);signal cellin_17_6 : std_logic_vector(1 downto 0);signal cellin_17_7 : std_logic_vector(1 downto 0);signal cellin_17_8 : std_logic_vector(0 downto 0);signal cellin_17_9 : std_logic_vector(0 downto 0);signal cellin_17_10 : std_logic_vector(0 downto 0);signal cellin_17_11 : std_logic_vector(0 downto 0);signal cellout_1_1 : std_logic_vector(3 downto 0);signal cellout_1_2 : std_logic_vector(3 downto 0);signal cellout_1_3 : std_logic_vector(3 downto 0);signal cellout_1_4 : std_logic_vector(3 downto 0);signal cellout_1_5 : std_logic_vector(2 downto 0);signal cellout_1_6 : std_logic_vector(3 downto 0);signal cellout_1_7 : std_logic_vector(2 downto 0);signal cellout_1_8 : std_logic_vector(0 downto 0);signal cellout_1_9 : std_logic_vector(1 downto 0);signal cellout_1_10 : std_logic_vector(0 downto 0);signal cellout_2_1 : std_logic_vector(2 downto 0);signal cellout_2_2 : std_logic_vector(2 downto 0);signal cellout_2_3 : std_logic_vector(2 downto 0);signal cellout_2_4 : std_logic_vector(2 downto 0);signal cellout_2_5 : std_logic_vector(1 downto 0);signal cellout_2_6 : std_logic_vector(2 downto 0);signal cellout_2_7 : std_logic_vector(0 downto 0);signal cellout_2_8 : std_logic_vector(0 downto 0);signal cellout_2_9 : std_logic_vector(1 downto 0);signal cellout_2_10 : std_logic_vector(0 downto 0);signal cellout_3_1 : std_logic_vector(1 downto 0);signal cellout_3_2 : std_logic_vector(1 downto 0);signal cellout_3_3 : std_logic_vector(1 downto 0);signal cellout_3_4 : std_logic_vector(1 downto 0);signal cellout_3_5 : std_logic_vector(1 downto 0);signal cellout_3_6 : std_logic_vector(0 downto 0);signal cellout_3_7 : std_logic_vector(0 downto 0);signal cellout_3_8 : std_logic_vector(0 downto 0);signal cellout_3_9 : std_logic_vector(1 downto 0);signal cellout_3_10 : std_logic_vector(0 downto 0);signal cellout_4_1 : std_logic_vector(1 downto 0);signal cellout_4_2 : std_logic_vector(1 downto 0);signal cellout_4_3 : std_logic_vector(1 downto 0);signal cellout_4_4 : std_logic_vector(1 downto 0);signal cellout_4_5 : std_logic_vector(1 downto 0);signal cellout_4_6 : std_logic_vector(0 downto 0);signal cellout_4_7 : std_logic_vector(0 downto 0);signal cellout_4_8 : std_logic_vector(0 downto 0);signal cellout_4_9 : std_logic_vector(1 downto 0);signal cellout_4_10 : std_logic_vector(0 downto 0);signal cellout_5_1 : std_logic_vector(1 downto 0);signal cellout_5_2 : std_logic_vector(1 downto 0);signal cellout_5_3 : std_logic_vector(2 downto 0);signal cellout_5_4 : std_logic_vector(1 downto 0);signal cellout_5_5 : std_logic_vector(1 downto 0);signal cellout_5_6 : std_logic_vector(1 downto 0);signal cellout_5_7 : std_logic_vector(1 downto 0);signal cellout_5_8 : std_logic_vector(1 downto 0);signal cellout_5_9 : std_logic_vector(1 downto 0);signal cellout_5_10 : std_logic_vector(1 downto 0);signal cellout_5_11 : std_logic_vector(0 downto 0);signal cellout_6_1 : std_logic_vector(1 downto 0);signal cellout_6_2 : std_logic_vector(1 downto 0);signal cellout_6_3 : std_logic_vector(0 downto 0);signal cellout_6_4 : std_logic_vector(1 downto 0);signal cellout_6_5 : std_logic_vector(1 downto 0);signal cellout_6_6 : std_logic_vector(1 downto 0);signal cellout_6_7 : std_logic_vector(1 downto 0);signal cellout_6_8 : std_logic_vector(1 downto 0);signal cellout_6_9 : std_logic_vector(1 downto 0);signal cellout_6_10 : std_logic_vector(1 downto 0);signal cellout_6_11 : std_logic_vector(0 downto 0);signal cellout_7_1 : std_logic_vector(1 downto 0);signal cellout_7_2 : std_logic_vector(1 downto 0);signal cellout_7_3 : std_logic_vector(1 downto 0);signal cellout_7_4 : std_logic_vector(1 downto 0);signal cellout_7_5 : std_logic_vector(1 downto 0);signal cellout_7_6 : std_logic_vector(1 downto 0);signal cellout_7_7 : std_logic_vector(1 downto 0);signal cellout_7_8 : std_logic_vector(0 downto 0);signal cellout_7_9 : std_logic_vector(1 downto 0);signal cellout_7_10 : std_logic_vector(1 downto 0);signal cellout_7_11 : std_logic_vector(0 downto 0);signal cellout_8_1 : std_logic_vector(1 downto 0);signal cellout_8_2 : std_logic_vector(1 downto 0);signal cellout_8_3 : std_logic_vector(1 downto 0);signal cellout_8_4 : std_logic_vector(1 downto 0);signal cellout_8_5 : std_logic_vector(1 downto 0);signal cellout_8_6 : std_logic_vector(1 downto 0);signal cellout_8_7 : std_logic_vector(1 downto 0);signal cellout_8_8 : std_logic_vector(0 downto 0);signal cellout_8_9 : std_logic_vector(1 downto 0);signal cellout_8_10 : std_logic_vector(1 downto 0);signal cellout_8_11 : std_logic_vector(0 downto 0);signal cellout_9_1 : std_logic_vector(1 downto 0);signal cellout_9_2 : std_logic_vector(1 downto 0);signal cellout_9_3 : std_logic_vector(2 downto 0);signal cellout_9_4 : std_logic_vector(1 downto 0);signal cellout_9_5 : std_logic_vector(1 downto 0);signal cellout_9_6 : std_logic_vector(2 downto 0);signal cellout_9_7 : std_logic_vector(2 downto 0);signal cellout_9_8 : std_logic_vector(1 downto 0);signal cellout_9_9 : std_logic_vector(2 downto 0);signal cellout_9_10 : std_logic_vector(0 downto 0);signal cellout_9_11 : std_logic_vector(1 downto 0);signal cellout_10_1 : std_logic_vector(1 downto 0);signal cellout_10_2 : std_logic_vector(1 downto 0);signal cellout_10_3 : std_logic_vector(1 downto 0);signal cellout_10_4 : std_logic_vector(1 downto 0);signal cellout_10_5 : std_logic_vector(1 downto 0);signal cellout_10_6 : std_logic_vector(1 downto 0);signal cellout_10_7 : std_logic_vector(1 downto 0);signal cellout_10_8 : std_logic_vector(1 downto 0);signal cellout_10_9 : std_logic_vector(0 downto 0);signal cellout_10_10 : std_logic_vector(0 downto 0);signal cellout_10_11 : std_logic_vector(1 downto 0);signal cellout_11_1 : std_logic_vector(1 downto 0);signal cellout_11_2 : std_logic_vector(1 downto 0);signal cellout_11_3 : std_logic_vector(1 downto 0);signal cellout_11_4 : std_logic_vector(1 downto 0);signal cellout_11_5 : std_logic_vector(1 downto 0);signal cellout_11_6 : std_logic_vector(1 downto 0);signal cellout_11_7 : std_logic_vector(1 downto 0);signal cellout_11_8 : std_logic_vector(1 downto 0);signal cellout_11_9 : std_logic_vector(0 downto 0);signal cellout_11_10 : std_logic_vector(0 downto 0);signal cellout_11_11 : std_logic_vector(1 downto 0);signal cellout_12_1 : std_logic_vector(2 downto 0);signal cellout_12_2 : std_logic_vector(2 downto 0);signal cellout_12_3 : std_logic_vector(1 downto 0);signal cellout_12_4 : std_logic_vector(1 downto 0);signal cellout_12_5 : std_logic_vector(2 downto 0);signal cellout_12_6 : std_logic_vector(1 downto 0);signal cellout_12_7 : std_logic_vector(1 downto 0);signal cellout_12_8 : std_logic_vector(1 downto 0);signal cellout_12_9 : std_logic_vector(0 downto 0);signal cellout_12_10 : std_logic_vector(0 downto 0);signal cellout_12_11 : std_logic_vector(1 downto 0);signal cellout_13_1 : std_logic_vector(5 downto 0);signal cellout_13_2 : std_logic_vector(5 downto 0);signal cellout_13_3 : std_logic_vector(5 downto 0);signal cellout_13_4 : std_logic_vector(5 downto 0);signal cellout_13_5 : std_logic_vector(4 downto 0);signal cellout_13_6 : std_logic_vector(4 downto 0);signal cellout_13_7 : std_logic_vector(2 downto 0);signal cellout_13_8 : std_logic_vector(3 downto 0);signal cellout_13_9 : std_logic_vector(0 downto 0);signal cellout_13_10 : std_logic_vector(2 downto 0);signal cellout_13_11 : std_logic_vector(0 downto 0);signal cellout_14_1 : std_logic_vector(3 downto 0);signal cellout_14_2 : std_logic_vector(3 downto 0);signal cellout_14_3 : std_logic_vector(3 downto 0);signal cellout_14_4 : std_logic_vector(2 downto 0);signal cellout_14_5 : std_logic_vector(3 downto 0);signal cellout_14_6 : std_logic_vector(3 downto 0);signal cellout_14_7 : std_logic_vector(1 downto 0);signal cellout_14_8 : std_logic_vector(1 downto 0);signal cellout_14_9 : std_logic_vector(1 downto 0);signal cellout_14_10 : std_logic_vector(0 downto 0);signal cellout_14_11 : std_logic_vector(0 downto 0);signal cellout_15_1 : std_logic_vector(2 downto 0);signal cellout_15_2 : std_logic_vector(2 downto 0);signal cellout_15_3 : std_logic_vector(2 downto 0);signal cellout_15_4 : std_logic_vector(1 downto 0);signal cellout_15_5 : std_logic_vector(2 downto 0);signal cellout_15_6 : std_logic_vector(1 downto 0);signal cellout_15_7 : std_logic_vector(1 downto 0);signal cellout_15_8 : std_logic_vector(2 downto 0);signal cellout_15_9 : std_logic_vector(0 downto 0);signal cellout_15_10 : std_logic_vector(0 downto 0);signal cellout_15_11 : std_logic_vector(0 downto 0);signal cellout_16_1 : std_logic_vector(1 downto 0);signal cellout_16_2 : std_logic_vector(1 downto 0);signal cellout_16_3 : std_logic_vector(1 downto 0);signal cellout_16_4 : std_logic_vector(1 downto 0);signal cellout_16_5 : std_logic_vector(1 downto 0);signal cellout_16_6 : std_logic_vector(1 downto 0);signal cellout_16_7 : std_logic_vector(1 downto 0);signal cellout_16_8 : std_logic_vector(0 downto 0);signal cellout_16_9 : std_logic_vector(0 downto 0);signal cellout_16_10 : std_logic_vector(0 downto 0);signal cellout_16_11 : std_logic_vector(0 downto 0);begincellin_1_10(0) <= in_1_10(0);cellin_1_9(0) <= in_1_9(0);cellin_1_9(1) <= in_1_9(1);cellin_1_8(0) <= in_1_8(0);cellin_1_8(1) <= in_1_8(1);cellin_1_8(2) <= in_1_8(2);cellin_1_7(0) <= in_1_7(0);cellin_1_7(1) <= in_1_7(1);cellin_1_7(2) <= in_1_7(2);cellin_1_7(3) <= in_1_7(3);cellin_1_6(0) <= in_1_6(0);cellin_1_6(1) <= in_1_6(1);cellin_1_6(2) <= in_1_6(2);cellin_1_6(3) <= in_1_6(3);cellin_1_6(4) <= in_1_6(4);cellin_1_5(0) <= in_1_5(0);cellin_1_5(1) <= in_1_5(1);cellin_1_5(2) <= in_1_5(2);cellin_1_5(3) <= in_1_5(3);cellin_1_5(4) <= in_1_5(4);cellin_1_5(5) <= in_1_5(5);cellin_1_4(0) <= in_1_4(0);cellin_1_4(1) <= in_1_4(1);cellin_1_4(2) <= in_1_4(2);cellin_1_4(3) <= in_1_4(3);cellin_1_4(4) <= in_1_4(4);cellin_1_4(5) <= in_1_4(5);cellin_1_3(0) <= in_1_3(0);cellin_1_3(1) <= in_1_3(1);cellin_1_3(2) <= in_1_3(2);cellin_1_3(3) <= in_1_3(3);cellin_1_3(4) <= in_1_3(4);cellin_1_3(5) <= in_1_3(5);cellin_1_2(0) <= in_1_2(0);cellin_1_2(1) <= in_1_2(1);cellin_1_2(2) <= in_1_2(2);cellin_1_2(3) <= in_1_2(3);cellin_1_2(4) <= in_1_2(4);cellin_1_2(5) <= in_1_2(5);cellin_1_1(0) <= in_1_1(0);cellin_1_1(1) <= in_1_1(1);cellin_1_1(2) <= in_1_1(2);cellin_1_1(3) <= in_1_1(3);cellin_1_1(4) <= in_1_1(4);cellin_1_1(5) <= in_1_1(5);cellin_5_11(0) <= in_5_11(0);cellin_5_10(0) <= in_5_10(0);cellin_5_9(0) <= in_5_9(0);cellin_5_9(1) <= in_5_9(1);cellin_5_8(0) <= in_5_8(0);cellin_5_8(1) <= in_5_8(1);cellin_5_7(0) <= in_5_7(0);cellin_5_7(1) <= in_5_7(1);cellin_5_6(0) <= in_5_6(0);cellin_5_6(1) <= in_5_6(1);cellin_5_5(0) <= in_5_5(0);cellin_5_4(0) <= in_5_4(0);cellin_7_8(0) <= in_7_8(0);cellin_7_7(0) <= in_7_7(0);cellin_7_6(0) <= in_7_6(0);cellin_7_5(0) <= in_7_5(0);cellin_7_4(0) <= in_7_4(0);cellin_7_3(0) <= in_7_3(0);cellin_9_11(0) <= in_9_11(0);cellin_9_10(0) <= in_9_10(0);cellin_9_9(0) <= in_9_9(0);cellin_9_9(1) <= in_9_9(1);cellin_9_8(0) <= in_9_8(0);cellin_9_8(1) <= in_9_8(1);cellin_9_7(0) <= in_9_7(0);cellin_9_7(1) <= in_9_7(1);cellin_9_6(0) <= in_9_6(0);cellin_9_6(1) <= in_9_6(1);cellin_9_5(0) <= in_9_5(0);cellin_9_4(0) <= in_9_4(0);cellin_13_10(0) <= in_13_10(0);cellin_13_9(0) <= in_13_9(0);cellin_13_9(1) <= in_13_9(1);cellin_13_8(0) <= in_13_8(0);cellin_13_8(1) <= in_13_8(1);cellin_13_8(2) <= in_13_8(2);cellin_13_7(0) <= in_13_7(0);cellin_13_7(1) <= in_13_7(1);cellin_13_7(2) <= in_13_7(2);cellin_13_7(3) <= in_13_7(3);cellin_13_6(0) <= in_13_6(0);cellin_13_6(1) <= in_13_6(1);cellin_13_6(2) <= in_13_6(2);cellin_13_6(3) <= in_13_6(3);cellin_13_6(4) <= in_13_6(4);cellin_13_5(0) <= in_13_5(0);cellin_13_5(1) <= in_13_5(1);cellin_13_5(2) <= in_13_5(2);cellin_13_5(3) <= in_13_5(3);cellin_13_5(4) <= in_13_5(4);cellin_13_5(5) <= in_13_5(5);cellin_13_4(0) <= in_13_4(0);cellin_13_4(1) <= in_13_4(1);cellin_13_4(2) <= in_13_4(2);cellin_13_4(3) <= in_13_4(3);cellin_13_4(4) <= in_13_4(4);cellin_13_4(5) <= in_13_4(5);cellin_13_3(0) <= in_13_3(0);cellin_13_3(1) <= in_13_3(1);cellin_13_3(2) <= in_13_3(2);cellin_13_3(3) <= in_13_3(3);cellin_13_3(4) <= in_13_3(4);cellin_13_3(5) <= in_13_3(5);cellin_13_2(0) <= in_13_2(0);cellin_13_2(1) <= in_13_2(1);cellin_13_2(2) <= in_13_2(2);cellin_13_2(3) <= in_13_2(3);cellin_13_2(4) <= in_13_2(4);cellin_13_2(5) <= in_13_2(5);cellin_13_1(0) <= in_13_1(0);cellin_13_1(1) <= in_13_1(1);cellin_13_1(2) <= in_13_1(2);cellin_13_1(3) <= in_13_1(3);cellin_13_1(4) <= in_13_1(4);cellin_13_1(5) <= in_13_1(5);cellin_1_5(6) <= '1';cellin_1_2(6) <= '1';cellin_1_1(6) <= '1';add_1_8_2_1_0: fa port map(cellin_1_8(2), cellin_1_8(1), cellin_1_8(0), cellout_1_8(0), cellout_1_7(0));add_1_7_3_2_1: fa port map(cellin_1_7(3), cellin_1_7(2), cellin_1_7(1), cellout_1_7(1), cellout_1_6(0));add_1_6_4_3_2: fa port map(cellin_1_6(4), cellin_1_6(3), cellin_1_6(2), cellout_1_6(1), cellout_1_5(0));add_1_5_5_4_3: fa port map(cellin_1_5(5), cellin_1_5(4), cellin_1_5(3), cellout_1_5(1), cellout_1_4(0));add_1_5_2_1_0: fa port map(cellin_1_5(2), cellin_1_5(1), cellin_1_5(0), cellout_1_5(2), cellout_1_4(1));add_1_4_5_4_3: fa port map(cellin_1_4(5), cellin_1_4(4), cellin_1_4(3), cellout_1_4(2), cellout_1_3(0));add_1_4_2_1_0: fa port map(cellin_1_4(2), cellin_1_4(1), cellin_1_4(0), cellout_1_4(3), cellout_1_3(1));add_1_3_5_4_3: fa port map(cellin_1_3(5), cellin_1_3(4), cellin_1_3(3), cellout_1_3(2), cellout_1_2(0));add_1_3_2_1_0: fa port map(cellin_1_3(2), cellin_1_3(1), cellin_1_3(0), cellout_1_3(3), cellout_1_2(1));add_1_2_5_4_3: fa port map(cellin_1_2(5), cellin_1_2(4), cellin_1_2(3), cellout_1_2(2), cellout_1_1(0));add_1_2_2_1_0: fa port map(cellin_1_2(2), cellin_1_2(1), cellin_1_2(0), cellout_1_2(3), cellout_1_1(1));add_1_1_5_4_3: fa_noc port map(cellin_1_1(5), cellin_1_1(4), cellin_1_1(3), cellout_1_1(2));add_1_1_2_1_0: fa_noc port map(cellin_1_1(2), cellin_1_1(1), cellin_1_1(0), cellout_1_1(3));add_2_7_2_1_0: fa port map(cellin_2_7(2), cellin_2_7(1), cellin_2_7(0), cellout_2_7(0), cellout_2_6(0));add_2_6_3_2_1: fa port map(cellin_2_6(3), cellin_2_6(2), cellin_2_6(1), cellout_2_6(1), cellout_2_5(0));add_2_5_2_1_0: fa port map(cellin_2_5(2), cellin_2_5(1), cellin_2_5(0), cellout_2_5(1), cellout_2_4(0));add_2_4_3_2_1: fa port map(cellin_2_4(3), cellin_2_4(2), cellin_2_4(1), cellout_2_4(1), cellout_2_3(0));add_2_3_3_2_1: fa port map(cellin_2_3(3), cellin_2_3(2), cellin_2_3(1), cellout_2_3(1), cellout_2_2(0));add_2_2_3_2_1: fa port map(cellin_2_2(3), cellin_2_2(2), cellin_2_2(1), cellout_2_2(1), cellout_2_1(0));add_2_1_3_2_1: fa_noc port map(cellin_2_1(3), cellin_2_1(2), cellin_2_1(1), cellout_2_1(1));add_3_6_2_1_0: fa port map(cellin_3_6(2), cellin_3_6(1), cellin_3_6(0), cellout_3_6(0), cellout_3_5(0));add_3_4_2_1_0: fa port map(cellin_3_4(2), cellin_3_4(1), cellin_3_4(0), cellout_3_4(1), cellout_3_3(0));add_3_3_2_1_0: fa port map(cellin_3_3(2), cellin_3_3(1), cellin_3_3(0), cellout_3_3(1), cellout_3_2(0));add_3_2_2_1_0: fa port map(cellin_3_2(2), cellin_3_2(1), cellin_3_2(0), cellout_3_2(1), cellout_3_1(0));add_3_1_2_1_0: fa_noc port map(cellin_3_1(2), cellin_3_1(1), cellin_3_1(0), cellout_3_1(1));add_5_9_3_2_1: fa port map(cellin_5_9(3), cellin_5_9(2), cellin_5_9(1), cellout_5_9(0), cellout_5_8(0));add_5_8_2_1_0: fa port map(cellin_5_8(2), cellin_5_8(1), cellin_5_8(0), cellout_5_8(1), cellout_5_7(0));add_5_7_2_1_0: fa port map(cellin_5_7(2), cellin_5_7(1), cellin_5_7(0), cellout_5_7(1), cellout_5_6(0));add_5_6_2_1_0: fa port map(cellin_5_6(2), cellin_5_6(1), cellin_5_6(0), cellout_5_6(1), cellout_5_5(0));add_5_5_2_1_0: fa port map(cellin_5_5(2), cellin_5_5(1), cellin_5_5(0), cellout_5_5(1), cellout_5_4(0));add_5_4_2_1_0: fa port map(cellin_5_4(2), cellin_5_4(1), cellin_5_4(0), cellout_5_4(1), cellout_5_3(0));add_6_3_2_1_0: fa port map(cellin_6_3(2), cellin_6_3(1), cellin_6_3(0), cellout_6_3(0), cellout_6_2(0));add_7_8_2_1_0: fa port map(cellin_7_8(2), cellin_7_8(1), cellin_7_8(0), cellout_7_8(0), cellout_7_7(0));add_7_7_2_1_0: fa port map(cellin_7_7(2), cellin_7_7(1), cellin_7_7(0), cellout_7_7(1), cellout_7_6(0));add_7_6_2_1_0: fa port map(cellin_7_6(2), cellin_7_6(1), cellin_7_6(0), cellout_7_6(1), cellout_7_5(0));add_7_5_2_1_0: fa port map(cellin_7_5(2), cellin_7_5(1), cellin_7_5(0), cellout_7_5(1), cellout_7_4(0));add_7_4_2_1_0: fa port map(cellin_7_4(2), cellin_7_4(1), cellin_7_4(0), cellout_7_4(1), cellout_7_3(0));add_9_10_2_1_0: fa port map(cellin_9_10(2), cellin_9_10(1), cellin_9_10(0), cellout_9_10(0), cellout_9_9(0));add_9_9_3_2_1: fa port map(cellin_9_9(3), cellin_9_9(2), cellin_9_9(1), cellout_9_9(1), cellout_9_8(0));add_9_8_2_1_0: fa port map(cellin_9_8(2), cellin_9_8(1), cellin_9_8(0), cellout_9_8(1), cellout_9_7(0));add_9_7_3_2_1: fa port map(cellin_9_7(3), cellin_9_7(2), cellin_9_7(1), cellout_9_7(1), cellout_9_6(0));add_9_6_3_2_1: fa port map(cellin_9_6(3), cellin_9_6(2), cellin_9_6(1), cellout_9_6(1), cellout_9_5(0));add_9_5_2_1_0: fa port map(cellin_9_5(2), cellin_9_5(1), cellin_9_5(0), cellout_9_5(1), cellout_9_4(0));add_9_4_2_1_0: fa port map(cellin_9_4(2), cellin_9_4(1), cellin_9_4(0), cellout_9_4(1), cellout_9_3(0));add_10_9_2_1_0: fa port map(cellin_10_9(2), cellin_10_9(1), cellin_10_9(0), cellout_10_9(0), cellout_10_8(0));add_10_7_2_1_0: fa port map(cellin_10_7(2), cellin_10_7(1), cellin_10_7(0), cellout_10_7(1), cellout_10_6(0));add_10_6_2_1_0: fa port map(cellin_10_6(2), cellin_10_6(1), cellin_10_6(0), cellout_10_6(1), cellout_10_5(0));add_10_3_2_1_0: fa port map(cellin_10_3(2), cellin_10_3(1), cellin_10_3(0), cellout_10_3(1), cellout_10_2(0));add_13_9_2_1_0: fa port map(cellin_13_9(2), cellin_13_9(1), cellin_13_9(0), cellout_13_9(0), cellout_13_8(0));add_13_8_4_3_2: fa port map(cellin_13_8(4), cellin_13_8(3), cellin_13_8(2), cellout_13_8(1), cellout_13_7(0));add_13_7_5_4_3: fa port map(cellin_13_7(5), cellin_13_7(4), cellin_13_7(3), cellout_13_7(1), cellout_13_6(0));add_13_7_2_1_0: fa port map(cellin_13_7(2), cellin_13_7(1), cellin_13_7(0), cellout_13_7(2), cellout_13_6(1));add_13_6_6_5_4: fa port map(cellin_13_6(6), cellin_13_6(5), cellin_13_6(4), cellout_13_6(2), cellout_13_5(0));add_13_6_3_2_1: fa port map(cellin_13_6(3), cellin_13_6(2), cellin_13_6(1), cellout_13_6(3), cellout_13_5(1));add_13_5_8_7_6: fa port map(cellin_13_5(8), cellin_13_5(7), cellin_13_5(6), cellout_13_5(2), cellout_13_4(0));add_13_5_5_4_3: fa port map(cellin_13_5(5), cellin_13_5(4), cellin_13_5(3), cellout_13_5(3), cellout_13_4(1));add_13_5_2_1_0: fa port map(cellin_13_5(2), cellin_13_5(1), cellin_13_5(0), cellout_13_5(4), cellout_13_4(2));add_13_4_7_6_5: fa port map(cellin_13_4(7), cellin_13_4(6), cellin_13_4(5), cellout_13_4(3), cellout_13_3(0));add_13_4_4_3_2: fa port map(cellin_13_4(4), cellin_13_4(3), cellin_13_4(2), cellout_13_4(4), cellout_13_3(1));add_13_3_7_6_5: fa port map(cellin_13_3(7), cellin_13_3(6), cellin_13_3(5), cellout_13_3(3), cellout_13_2(0));add_13_3_4_3_2: fa port map(cellin_13_3(4), cellin_13_3(3), cellin_13_3(2), cellout_13_3(4), cellout_13_2(1));add_13_2_8_7_6: fa port map(cellin_13_2(8), cellin_13_2(7), cellin_13_2(6), cellout_13_2(3), cellout_13_1(0));add_13_2_5_4_3: fa port map(cellin_13_2(5), cellin_13_2(4), cellin_13_2(3), cellout_13_2(4), cellout_13_1(1));add_13_2_2_1_0: fa port map(cellin_13_2(2), cellin_13_2(1), cellin_13_2(0), cellout_13_2(5), cellout_13_1(2));add_13_1_8_7_6: fa_noc port map(cellin_13_1(8), cellin_13_1(7), cellin_13_1(6), cellout_13_1(3));add_13_1_5_4_3: fa_noc port map(cellin_13_1(5), cellin_13_1(4), cellin_13_1(3), cellout_13_1(4));add_13_1_2_1_0: fa_noc port map(cellin_13_1(2), cellin_13_1(1), cellin_13_1(0), cellout_13_1(5));add_14_10_2_1_0: fa port map(cellin_14_10(2), cellin_14_10(1), cellin_14_10(0), cellout_14_10(0), cellout_14_9(0));add_14_8_3_2_1: fa port map(cellin_14_8(3), cellin_14_8(2), cellin_14_8(1), cellout_14_8(0), cellout_14_7(0));add_14_7_2_1_0: fa port map(cellin_14_7(2), cellin_14_7(1), cellin_14_7(0), cellout_14_7(1), cellout_14_6(0));add_14_6_4_3_2: fa port map(cellin_14_6(4), cellin_14_6(3), cellin_14_6(2), cellout_14_6(1), cellout_14_5(0));add_14_5_4_3_2: fa port map(cellin_14_5(4), cellin_14_5(3), cellin_14_5(2), cellout_14_5(1), cellout_14_4(0));add_14_4_5_4_3: fa port map(cellin_14_4(5), cellin_14_4(4), cellin_14_4(3), cellout_14_4(1), cellout_14_3(0));add_14_4_2_1_0: fa port map(cellin_14_4(2), cellin_14_4(1), cellin_14_4(0), cellout_14_4(2), cellout_14_3(1));add_14_3_5_4_3: fa port map(cellin_14_3(5), cellin_14_3(4), cellin_14_3(3), cellout_14_3(2), cellout_14_2(0));add_14_3_2_1_0: fa port map(cellin_14_3(2), cellin_14_3(1), cellin_14_3(0), cellout_14_3(3), cellout_14_2(1));add_14_2_5_4_3: fa port map(cellin_14_2(5), cellin_14_2(4), cellin_14_2(3), cellout_14_2(2), cellout_14_1(0));add_14_2_2_1_0: fa port map(cellin_14_2(2), cellin_14_2(1), cellin_14_2(0), cellout_14_2(3), cellout_14_1(1));add_14_1_5_4_3: fa_noc port map(cellin_14_1(5), cellin_14_1(4), cellin_14_1(3), cellout_14_1(2));add_14_1_2_1_0: fa_noc port map(cellin_14_1(2), cellin_14_1(1), cellin_14_1(0), cellout_14_1(3));add_15_6_3_2_1: fa port map(cellin_15_6(3), cellin_15_6(2), cellin_15_6(1), cellout_15_6(0), cellout_15_5(0));add_15_5_3_2_1: fa port map(cellin_15_5(3), cellin_15_5(2), cellin_15_5(1), cellout_15_5(1), cellout_15_4(0));add_15_4_2_1_0: fa port map(cellin_15_4(2), cellin_15_4(1), cellin_15_4(0), cellout_15_4(1), cellout_15_3(0));add_15_3_3_2_1: fa port map(cellin_15_3(3), cellin_15_3(2), cellin_15_3(1), cellout_15_3(1), cellout_15_2(0));add_15_2_3_2_1: fa port map(cellin_15_2(3), cellin_15_2(2), cellin_15_2(1), cellout_15_2(1), cellout_15_1(0));add_15_1_3_2_1: fa_noc port map(cellin_15_1(3), cellin_15_1(2), cellin_15_1(1), cellout_15_1(1));add_16_8_2_1_0: fa port map(cellin_16_8(2), cellin_16_8(1), cellin_16_8(0), cellout_16_8(0), cellout_16_7(0));add_16_5_2_1_0: fa port map(cellin_16_5(2), cellin_16_5(1), cellin_16_5(0), cellout_16_5(1), cellout_16_4(0));add_16_3_2_1_0: fa port map(cellin_16_3(2), cellin_16_3(1), cellin_16_3(0), cellout_16_3(1), cellout_16_2(0));add_16_2_2_1_0: fa port map(cellin_16_2(2), cellin_16_2(1), cellin_16_2(0), cellout_16_2(1), cellout_16_1(0));add_16_1_2_1_0: fa_noc port map(cellin_16_1(2), cellin_16_1(1), cellin_16_1(0), cellout_16_1(1));add_3_5_1_0: ha port map(cellin_3_5(1), cellin_3_5(0), cellout_3_5(1), cellout_3_4(0));add_6_2_1_0: ha port map(cellin_6_2(1), cellin_6_2(0), cellout_6_2(1), cellout_6_1(0));add_6_1_1_0: ha_noc port map(cellin_6_1(1), cellin_6_1(0), cellout_6_1(1));add_7_3_1_0: ha port map(cellin_7_3(1), cellin_7_3(0), cellout_7_3(1), cellout_7_2(0));add_7_2_1_0: ha port map(cellin_7_2(1), cellin_7_2(0), cellout_7_2(1), cellout_7_1(0));add_7_1_1_0: ha_noc port map(cellin_7_1(1), cellin_7_1(0), cellout_7_1(1));add_10_8_1_0: ha port map(cellin_10_8(1), cellin_10_8(0), cellout_10_8(1), cellout_10_7(0));add_10_5_1_0: ha port map(cellin_10_5(1), cellin_10_5(0), cellout_10_5(1), cellout_10_4(0));add_10_4_1_0: ha port map(cellin_10_4(1), cellin_10_4(0), cellout_10_4(1), cellout_10_3(0));add_10_2_1_0: ha port map(cellin_10_2(1), cellin_10_2(0), cellout_10_2(1), cellout_10_1(0));add_10_1_1_0: ha_noc port map(cellin_10_1(1), cellin_10_1(0), cellout_10_1(1));add_13_11_1_0: ha port map(cellin_13_11(1), cellin_13_11(0), cellout_13_11(0), cellout_13_10(0));add_13_4_1_0: ha port map(cellin_13_4(1), cellin_13_4(0), cellout_13_4(5), cellout_13_3(2));add_13_3_1_0: ha port map(cellin_13_3(1), cellin_13_3(0), cellout_13_3(5), cellout_13_2(2));add_15_9_1_0: ha port map(cellin_15_9(1), cellin_15_9(0), cellout_15_9(0), cellout_15_8(0));add_16_7_1_0: ha port map(cellin_16_7(1), cellin_16_7(0), cellout_16_7(1), cellout_16_6(0));add_16_6_1_0: ha port map(cellin_16_6(1), cellin_16_6(0), cellout_16_6(1), cellout_16_5(0));add_16_4_1_0: ha port map(cellin_16_4(1), cellin_16_4(0), cellout_16_4(1), cellout_16_3(0));cellout_1_10(0) <= cellin_1_10(0);cellout_1_9(0) <= cellin_1_9(1);cellout_1_9(1) <= cellin_1_9(0);cellout_1_7(2) <= cellin_1_7(0);cellout_1_6(2) <= cellin_1_6(1);cellout_1_6(3) <= cellin_1_6(0);cellout_2_10(0) <= cellin_2_10(0);cellout_2_9(0) <= cellin_2_9(1);cellout_2_9(1) <= cellin_2_9(0);cellout_2_8(0) <= cellin_2_8(0);cellout_2_6(2) <= cellin_2_6(0);cellout_2_4(2) <= cellin_2_4(0);cellout_2_3(2) <= cellin_2_3(0);cellout_2_2(2) <= cellin_2_2(0);cellout_2_1(2) <= cellin_2_1(0);cellout_3_10(0) <= cellin_3_10(0);cellout_3_9(0) <= cellin_3_9(1);cellout_3_9(1) <= cellin_3_9(0);cellout_3_8(0) <= cellin_3_8(0);cellout_3_7(0) <= cellin_3_7(0);cellout_4_10(0) <= cellin_4_10(0);cellout_4_9(0) <= cellin_4_9(1);cellout_4_9(1) <= cellin_4_9(0);cellout_4_8(0) <= cellin_4_8(0);cellout_4_7(0) <= cellin_4_7(0);cellout_4_6(0) <= cellin_4_6(0);cellout_4_5(0) <= cellin_4_5(1);cellout_4_5(1) <= cellin_4_5(0);cellout_4_4(0) <= cellin_4_4(1);cellout_4_4(1) <= cellin_4_4(0);cellout_4_3(0) <= cellin_4_3(1);cellout_4_3(1) <= cellin_4_3(0);cellout_4_2(0) <= cellin_4_2(1);cellout_4_2(1) <= cellin_4_2(0);cellout_4_1(0) <= cellin_4_1(1);cellout_4_1(1) <= cellin_4_1(0);cellout_5_11(0) <= cellin_5_11(0);cellout_5_10(0) <= cellin_5_10(1);cellout_5_10(1) <= cellin_5_10(0);cellout_5_9(1) <= cellin_5_9(0);cellout_5_3(1) <= cellin_5_3(1);cellout_5_3(2) <= cellin_5_3(0);cellout_5_2(0) <= cellin_5_2(1);cellout_5_2(1) <= cellin_5_2(0);cellout_5_1(0) <= cellin_5_1(1);cellout_5_1(1) <= cellin_5_1(0);cellout_6_11(0) <= cellin_6_11(0);cellout_6_10(0) <= cellin_6_10(1);cellout_6_10(1) <= cellin_6_10(0);cellout_6_9(0) <= cellin_6_9(1);cellout_6_9(1) <= cellin_6_9(0);cellout_6_8(0) <= cellin_6_8(1);cellout_6_8(1) <= cellin_6_8(0);cellout_6_7(0) <= cellin_6_7(1);cellout_6_7(1) <= cellin_6_7(0);cellout_6_6(0) <= cellin_6_6(1);cellout_6_6(1) <= cellin_6_6(0);cellout_6_5(0) <= cellin_6_5(1);cellout_6_5(1) <= cellin_6_5(0);cellout_6_4(0) <= cellin_6_4(1);cellout_6_4(1) <= cellin_6_4(0);cellout_7_11(0) <= cellin_7_11(0);cellout_7_10(0) <= cellin_7_10(1);cellout_7_10(1) <= cellin_7_10(0);cellout_7_9(0) <= cellin_7_9(1);cellout_7_9(1) <= cellin_7_9(0);cellout_8_11(0) <= cellin_8_11(0);cellout_8_10(0) <= cellin_8_10(1);cellout_8_10(1) <= cellin_8_10(0);cellout_8_9(0) <= cellin_8_9(1);cellout_8_9(1) <= cellin_8_9(0);cellout_8_8(0) <= cellin_8_8(0);cellout_8_7(0) <= cellin_8_7(1);cellout_8_7(1) <= cellin_8_7(0);cellout_8_6(0) <= cellin_8_6(1);cellout_8_6(1) <= cellin_8_6(0);cellout_8_5(0) <= cellin_8_5(1);cellout_8_5(1) <= cellin_8_5(0);cellout_8_4(0) <= cellin_8_4(1);cellout_8_4(1) <= cellin_8_4(0);cellout_8_3(0) <= cellin_8_3(1);cellout_8_3(1) <= cellin_8_3(0);cellout_8_2(0) <= cellin_8_2(1);cellout_8_2(1) <= cellin_8_2(0);cellout_8_1(0) <= cellin_8_1(1);cellout_8_1(1) <= cellin_8_1(0);cellout_9_11(0) <= cellin_9_11(1);cellout_9_11(1) <= cellin_9_11(0);cellout_9_9(2) <= cellin_9_9(0);cellout_9_7(2) <= cellin_9_7(0);cellout_9_6(2) <= cellin_9_6(0);cellout_9_3(1) <= cellin_9_3(1);cellout_9_3(2) <= cellin_9_3(0);cellout_9_2(0) <= cellin_9_2(1);cellout_9_2(1) <= cellin_9_2(0);cellout_9_1(0) <= cellin_9_1(1);cellout_9_1(1) <= cellin_9_1(0);cellout_10_11(0) <= cellin_10_11(1);cellout_10_11(1) <= cellin_10_11(0);cellout_10_10(0) <= cellin_10_10(0);cellout_11_11(0) <= cellin_11_11(1);cellout_11_11(1) <= cellin_11_11(0);cellout_11_10(0) <= cellin_11_10(0);cellout_11_9(0) <= cellin_11_9(0);cellout_11_8(0) <= cellin_11_8(1);cellout_11_8(1) <= cellin_11_8(0);cellout_11_7(0) <= cellin_11_7(1);cellout_11_7(1) <= cellin_11_7(0);cellout_11_6(0) <= cellin_11_6(1);cellout_11_6(1) <= cellin_11_6(0);cellout_11_5(0) <= cellin_11_5(1);cellout_11_5(1) <= cellin_11_5(0);cellout_11_4(0) <= cellin_11_4(1);cellout_11_4(1) <= cellin_11_4(0);cellout_11_3(0) <= cellin_11_3(1);cellout_11_3(1) <= cellin_11_3(0);cellout_11_2(0) <= cellin_11_2(1);cellout_11_2(1) <= cellin_11_2(0);cellout_11_1(0) <= cellin_11_1(1);cellout_11_1(1) <= cellin_11_1(0);cellout_12_11(0) <= cellin_12_11(1);cellout_12_11(1) <= cellin_12_11(0);cellout_12_10(0) <= cellin_12_10(0);cellout_12_9(0) <= cellin_12_9(0);cellout_12_8(0) <= cellin_12_8(1);cellout_12_8(1) <= cellin_12_8(0);cellout_12_7(0) <= cellin_12_7(1);cellout_12_7(1) <= cellin_12_7(0);cellout_12_6(0) <= cellin_12_6(1);cellout_12_6(1) <= cellin_12_6(0);cellout_12_5(0) <= cellin_12_5(1);cellout_12_5(1) <= cellin_12_5(0);cellout_12_4(0) <= cellin_12_4(1);cellout_12_4(1) <= cellin_12_4(0);cellout_12_3(0) <= cellin_12_3(1);cellout_12_3(1) <= cellin_12_3(0);cellout_12_2(0) <= cellin_12_2(1);cellout_12_2(1) <= cellin_12_2(0);cellout_12_1(0) <= cellin_12_1(1);cellout_12_1(1) <= cellin_12_1(0);cellout_13_10(1) <= cellin_13_10(1);cellout_13_10(2) <= cellin_13_10(0);cellout_13_8(2) <= cellin_13_8(1);cellout_13_8(3) <= cellin_13_8(0);cellout_13_6(4) <= cellin_13_6(0);cellout_14_11(0) <= cellin_14_11(0);cellout_14_9(1) <= cellin_14_9(0);cellout_14_8(1) <= cellin_14_8(0);cellout_14_6(2) <= cellin_14_6(1);cellout_14_6(3) <= cellin_14_6(0);cellout_14_5(2) <= cellin_14_5(1);cellout_14_5(3) <= cellin_14_5(0);cellout_15_11(0) <= cellin_15_11(0);cellout_15_10(0) <= cellin_15_10(0);cellout_15_8(1) <= cellin_15_8(1);cellout_15_8(2) <= cellin_15_8(0);cellout_15_7(0) <= cellin_15_7(1);cellout_15_7(1) <= cellin_15_7(0);cellout_15_6(1) <= cellin_15_6(0);cellout_15_5(2) <= cellin_15_5(0);cellout_15_3(2) <= cellin_15_3(0);cellout_15_2(2) <= cellin_15_2(0);cellout_15_1(2) <= cellin_15_1(0);cellout_16_11(0) <= cellin_16_11(0);cellout_16_10(0) <= cellin_16_10(0);cellout_16_9(0) <= cellin_16_9(0);reg_2_10_0: dff port map(clk, reset, cellout_2_10(0), cellin_3_10(0));reg_2_9_0: dff port map(clk, reset, cellout_2_9(0), cellin_3_9(0));reg_2_9_1: dff port map(clk, reset, cellout_2_9(1), cellin_3_9(1));reg_2_8_0: dff port map(clk, reset, cellout_2_8(0), cellin_3_8(0));reg_2_7_0: dff port map(clk, reset, cellout_2_7(0), cellin_3_7(0));reg_2_6_0: dff port map(clk, reset, cellout_2_6(0), cellin_3_6(0));reg_2_6_1: dff port map(clk, reset, cellout_2_6(1), cellin_3_6(1));reg_2_6_2: dff port map(clk, reset, cellout_2_6(2), cellin_3_6(2));reg_2_5_0: dff port map(clk, reset, cellout_2_5(0), cellin_3_5(0));reg_2_5_1: dff port map(clk, reset, cellout_2_5(1), cellin_3_5(1));reg_2_4_0: dff port map(clk, reset, cellout_2_4(0), cellin_3_4(0));reg_2_4_1: dff port map(clk, reset, cellout_2_4(1), cellin_3_4(1));reg_2_4_2: dff port map(clk, reset, cellout_2_4(2), cellin_3_4(2));reg_2_3_0: dff port map(clk, reset, cellout_2_3(0), cellin_3_3(0));reg_2_3_1: dff port map(clk, reset, cellout_2_3(1), cellin_3_3(1));reg_2_3_2: dff port map(clk, reset, cellout_2_3(2), cellin_3_3(2));reg_2_2_0: dff port map(clk, reset, cellout_2_2(0), cellin_3_2(0));reg_2_2_1: dff port map(clk, reset, cellout_2_2(1), cellin_3_2(1));reg_2_2_2: dff port map(clk, reset, cellout_2_2(2), cellin_3_2(2));reg_2_1_0: dff port map(clk, reset, cellout_2_1(0), cellin_3_1(0));reg_2_1_1: dff port map(clk, reset, cellout_2_1(1), cellin_3_1(1));reg_2_1_2: dff port map(clk, reset, cellout_2_1(2), cellin_3_1(2));reg_4_10_0: dff port map(clk, reset, cellout_4_10(0), cellin_5_10(1));reg_4_9_0: dff port map(clk, reset, cellout_4_9(0), cellin_5_9(2));reg_4_9_1: dff port map(clk, reset, cellout_4_9(1), cellin_5_9(3));reg_4_8_0: dff port map(clk, reset, cellout_4_8(0), cellin_5_8(2));reg_4_7_0: dff port map(clk, reset, cellout_4_7(0), cellin_5_7(2));reg_4_6_0: dff port map(clk, reset, cellout_4_6(0), cellin_5_6(2));reg_4_5_0: dff port map(clk, reset, cellout_4_5(0), cellin_5_5(1));reg_4_5_1: dff port map(clk, reset, cellout_4_5(1), cellin_5_5(2));reg_4_4_0: dff port map(clk, reset, cellout_4_4(0), cellin_5_4(1));reg_4_4_1: dff port map(clk, reset, cellout_4_4(1), cellin_5_4(2));reg_4_3_0: dff port map(clk, reset, cellout_4_3(0), cellin_5_3(0));reg_4_3_1: dff port map(clk, reset, cellout_4_3(1), cellin_5_3(1));reg_4_2_0: dff port map(clk, reset, cellout_4_2(0), cellin_5_2(0));reg_4_2_1: dff port map(clk, reset, cellout_4_2(1), cellin_5_2(1));reg_4_1_0: dff port map(clk, reset, cellout_4_1(0), cellin_5_1(0));reg_4_1_1: dff port map(clk, reset, cellout_4_1(1), cellin_5_1(1));reg_6_11_0: dff port map(clk, reset, cellout_6_11(0), cellin_7_11(0));reg_6_10_0: dff port map(clk, reset, cellout_6_10(0), cellin_7_10(0));reg_6_10_1: dff port map(clk, reset, cellout_6_10(1), cellin_7_10(1));reg_6_9_0: dff port map(clk, reset, cellout_6_9(0), cellin_7_9(0));reg_6_9_1: dff port map(clk, reset, cellout_6_9(1), cellin_7_9(1));reg_6_8_0: dff port map(clk, reset, cellout_6_8(0), cellin_7_8(1));reg_6_8_1: dff port map(clk, reset, cellout_6_8(1), cellin_7_8(2));reg_6_7_0: dff port map(clk, reset, cellout_6_7(0), cellin_7_7(1));reg_6_7_1: dff port map(clk, reset, cellout_6_7(1), cellin_7_7(2));reg_6_6_0: dff port map(clk, reset, cellout_6_6(0), cellin_7_6(1));reg_6_6_1: dff port map(clk, reset, cellout_6_6(1), cellin_7_6(2));reg_6_5_0: dff port map(clk, reset, cellout_6_5(0), cellin_7_5(1));reg_6_5_1: dff port map(clk, reset, cellout_6_5(1), cellin_7_5(2));reg_6_4_0: dff port map(clk, reset, cellout_6_4(0), cellin_7_4(1));reg_6_4_1: dff port map(clk, reset, cellout_6_4(1), cellin_7_4(2));reg_6_3_0: dff port map(clk, reset, cellout_6_3(0), cellin_7_3(1));reg_6_2_0: dff port map(clk, reset, cellout_6_2(0), cellin_7_2(0));reg_6_2_1: dff port map(clk, reset, cellout_6_2(1), cellin_7_2(1));reg_6_1_0: dff port map(clk, reset, cellout_6_1(0), cellin_7_1(0));reg_6_1_1: dff port map(clk, reset, cellout_6_1(1), cellin_7_1(1));reg_8_11_0: dff port map(clk, reset, cellout_8_11(0), cellin_9_11(1));reg_8_10_0: dff port map(clk, reset, cellout_8_10(0), cellin_9_10(1));reg_8_10_1: dff port map(clk, reset, cellout_8_10(1), cellin_9_10(2));reg_8_9_0: dff port map(clk, reset, cellout_8_9(0), cellin_9_9(2));reg_8_9_1: dff port map(clk, reset, cellout_8_9(1), cellin_9_9(3));reg_8_8_0: dff port map(clk, reset, cellout_8_8(0), cellin_9_8(2));reg_8_7_0: dff port map(clk, reset, cellout_8_7(0), cellin_9_7(2));reg_8_7_1: dff port map(clk, reset, cellout_8_7(1), cellin_9_7(3));reg_8_6_0: dff port map(clk, reset, cellout_8_6(0), cellin_9_6(2));reg_8_6_1: dff port map(clk, reset, cellout_8_6(1), cellin_9_6(3));reg_8_5_0: dff port map(clk, reset, cellout_8_5(0), cellin_9_5(1));reg_8_5_1: dff port map(clk, reset, cellout_8_5(1), cellin_9_5(2));reg_8_4_0: dff port map(clk, reset, cellout_8_4(0), cellin_9_4(1));reg_8_4_1: dff port map(clk, reset, cellout_8_4(1), cellin_9_4(2));reg_8_3_0: dff port map(clk, reset, cellout_8_3(0), cellin_9_3(0));reg_8_3_1: dff port map(clk, reset, cellout_8_3(1), cellin_9_3(1));reg_8_2_0: dff port map(clk, reset, cellout_8_2(0), cellin_9_2(0));reg_8_2_1: dff port map(clk, reset, cellout_8_2(1), cellin_9_2(1));reg_8_1_0: dff port map(clk, reset, cellout_8_1(0), cellin_9_1(0));reg_8_1_1: dff port map(clk, reset, cellout_8_1(1), cellin_9_1(1));reg_10_11_0: dff port map(clk, reset, cellout_10_11(0), cellin_11_11(0));reg_10_11_1: dff port map(clk, reset, cellout_10_11(1), cellin_11_11(1));reg_10_10_0: dff port map(clk, reset, cellout_10_10(0), cellin_11_10(0));reg_10_9_0: dff port map(clk, reset, cellout_10_9(0), cellin_11_9(0));reg_10_8_0: dff port map(clk, reset, cellout_10_8(0), cellin_11_8(0));reg_10_8_1: dff port map(clk, reset, cellout_10_8(1), cellin_11_8(1));reg_10_7_0: dff port map(clk, reset, cellout_10_7(0), cellin_11_7(0));reg_10_7_1: dff port map(clk, reset, cellout_10_7(1), cellin_11_7(1));reg_10_6_0: dff port map(clk, reset, cellout_10_6(0), cellin_11_6(0));reg_10_6_1: dff port map(clk, reset, cellout_10_6(1), cellin_11_6(1));reg_10_5_0: dff port map(clk, reset, cellout_10_5(0), cellin_11_5(0));reg_10_5_1: dff port map(clk, reset, cellout_10_5(1), cellin_11_5(1));reg_10_4_0: dff port map(clk, reset, cellout_10_4(0), cellin_11_4(0));reg_10_4_1: dff port map(clk, reset, cellout_10_4(1), cellin_11_4(1));reg_10_3_0: dff port map(clk, reset, cellout_10_3(0), cellin_11_3(0));reg_10_3_1: dff port map(clk, reset, cellout_10_3(1), cellin_11_3(1));reg_10_2_0: dff port map(clk, reset, cellout_10_2(0), cellin_11_2(0));reg_10_2_1: dff port map(clk, reset, cellout_10_2(1), cellin_11_2(1));reg_10_1_0: dff port map(clk, reset, cellout_10_1(0), cellin_11_1(0));reg_10_1_1: dff port map(clk, reset, cellout_10_1(1), cellin_11_1(1));reg_12_11_0: dff port map(clk, reset, cellout_12_11(0), cellin_13_11(0));reg_12_11_1: dff port map(clk, reset, cellout_12_11(1), cellin_13_11(1));reg_12_10_0: dff port map(clk, reset, cellout_12_10(0), cellin_13_10(1));reg_12_9_0: dff port map(clk, reset, cellout_12_9(0), cellin_13_9(2));reg_12_8_0: dff port map(clk, reset, cellout_12_8(0), cellin_13_8(3));reg_12_8_1: dff port map(clk, reset, cellout_12_8(1), cellin_13_8(4));reg_12_7_0: dff port map(clk, reset, cellout_12_7(0), cellin_13_7(4));reg_12_7_1: dff port map(clk, reset, cellout_12_7(1), cellin_13_7(5));reg_12_6_0: dff port map(clk, reset, cellout_12_6(0), cellin_13_6(5));reg_12_6_1: dff port map(clk, reset, cellout_12_6(1), cellin_13_6(6));reg_12_5_0: dff port map(clk, reset, cellout_12_5(0), cellin_13_5(6));reg_12_5_1: dff port map(clk, reset, cellout_12_5(1), cellin_13_5(7));reg_12_4_0: dff port map(clk, reset, cellout_12_4(0), cellin_13_4(6));reg_12_4_1: dff port map(clk, reset, cellout_12_4(1), cellin_13_4(7));reg_12_3_0: dff port map(clk, reset, cellout_12_3(0), cellin_13_3(6));reg_12_3_1: dff port map(clk, reset, cellout_12_3(1), cellin_13_3(7));reg_12_2_0: dff port map(clk, reset, cellout_12_2(0), cellin_13_2(6));reg_12_2_1: dff port map(clk, reset, cellout_12_2(1), cellin_13_2(7));reg_12_1_0: dff port map(clk, reset, cellout_12_1(0), cellin_13_1(6));reg_12_1_1: dff port map(clk, reset, cellout_12_1(1), cellin_13_1(7));reg_14_11_0: dff port map(clk, reset, cellout_14_11(0), cellin_15_11(0));reg_14_10_0: dff port map(clk, reset, cellout_14_10(0), cellin_15_10(0));reg_14_9_0: dff port map(clk, reset, cellout_14_9(0), cellin_15_9(0));reg_14_9_1: dff port map(clk, reset, cellout_14_9(1), cellin_15_9(1));reg_14_8_0: dff port map(clk, reset, cellout_14_8(0), cellin_15_8(0));reg_14_8_1: dff port map(clk, reset, cellout_14_8(1), cellin_15_8(1));reg_14_7_0: dff port map(clk, reset, cellout_14_7(0), cellin_15_7(0));reg_14_7_1: dff port map(clk, reset, cellout_14_7(1), cellin_15_7(1));reg_14_6_0: dff port map(clk, reset, cellout_14_6(0), cellin_15_6(0));reg_14_6_1: dff port map(clk, reset, cellout_14_6(1), cellin_15_6(1));reg_14_6_2: dff port map(clk, reset, cellout_14_6(2), cellin_15_6(2));reg_14_6_3: dff port map(clk, reset, cellout_14_6(3), cellin_15_6(3));reg_14_5_0: dff port map(clk, reset, cellout_14_5(0), cellin_15_5(0));reg_14_5_1: dff port map(clk, reset, cellout_14_5(1), cellin_15_5(1));reg_14_5_2: dff port map(clk, reset, cellout_14_5(2), cellin_15_5(2));reg_14_5_3: dff port map(clk, reset, cellout_14_5(3), cellin_15_5(3));reg_14_4_0: dff port map(clk, reset, cellout_14_4(0), cellin_15_4(0));reg_14_4_1: dff port map(clk, reset, cellout_14_4(1), cellin_15_4(1));reg_14_4_2: dff port map(clk, reset, cellout_14_4(2), cellin_15_4(2));reg_14_3_0: dff port map(clk, reset, cellout_14_3(0), cellin_15_3(0));reg_14_3_1: dff port map(clk, reset, cellout_14_3(1), cellin_15_3(1));reg_14_3_2: dff port map(clk, reset, cellout_14_3(2), cellin_15_3(2));reg_14_3_3: dff port map(clk, reset, cellout_14_3(3), cellin_15_3(3));reg_14_2_0: dff port map(clk, reset, cellout_14_2(0), cellin_15_2(0));reg_14_2_1: dff port map(clk, reset, cellout_14_2(1), cellin_15_2(1));reg_14_2_2: dff port map(clk, reset, cellout_14_2(2), cellin_15_2(2));reg_14_2_3: dff port map(clk, reset, cellout_14_2(3), cellin_15_2(3));reg_14_1_0: dff port map(clk, reset, cellout_14_1(0), cellin_15_1(0));reg_14_1_1: dff port map(clk, reset, cellout_14_1(1), cellin_15_1(1));reg_14_1_2: dff port map(clk, reset, cellout_14_1(2), cellin_15_1(2));reg_14_1_3: dff port map(clk, reset, cellout_14_1(3), cellin_15_1(3));reg_16_11_0: dff port map(clk, reset, cellout_16_11(0), cellin_17_11(0));reg_16_10_0: dff port map(clk, reset, cellout_16_10(0), cellin_17_10(0));reg_16_9_0: dff port map(clk, reset, cellout_16_9(0), cellin_17_9(0));reg_16_8_0: dff port map(clk, reset, cellout_16_8(0), cellin_17_8(0));reg_16_7_0: dff port map(clk, reset, cellout_16_7(0), cellin_17_7(0));reg_16_7_1: dff port map(clk, reset, cellout_16_7(1), cellin_17_7(1));reg_16_6_0: dff port map(clk, reset, cellout_16_6(0), cellin_17_6(0));reg_16_6_1: dff port map(clk, reset, cellout_16_6(1), cellin_17_6(1));reg_16_5_0: dff port map(clk, reset, cellout_16_5(0), cellin_17_5(0));reg_16_5_1: dff port map(clk, reset, cellout_16_5(1), cellin_17_5(1));reg_16_4_0: dff port map(clk, reset, cellout_16_4(0), cellin_17_4(0));reg_16_4_1: dff port map(clk, reset, cellout_16_4(1), cellin_17_4(1));reg_16_3_0: dff port map(clk, reset, cellout_16_3(0), cellin_17_3(0));reg_16_3_1: dff port map(clk, reset, cellout_16_3(1), cellin_17_3(1));reg_16_2_0: dff port map(clk, reset, cellout_16_2(0), cellin_17_2(0));reg_16_2_1: dff port map(clk, reset, cellout_16_2(1), cellin_17_2(1));reg_16_1_0: dff port map(clk, reset, cellout_16_1(0), cellin_17_1(0));reg_16_1_1: dff port map(clk, reset, cellout_16_1(1), cellin_17_1(1));cellin_2_10(0) <= cellout_1_10(0);cellin_2_9(0) <= cellout_1_9(0);cellin_2_9(1) <= cellout_1_9(1);cellin_2_8(0) <= cellout_1_8(0);cellin_2_7(0) <= cellout_1_7(0);cellin_2_7(1) <= cellout_1_7(1);cellin_2_7(2) <= cellout_1_7(2);cellin_2_6(0) <= cellout_1_6(0);cellin_2_6(1) <= cellout_1_6(1);cellin_2_6(2) <= cellout_1_6(2);cellin_2_6(3) <= cellout_1_6(3);cellin_2_5(0) <= cellout_1_5(0);cellin_2_5(1) <= cellout_1_5(1);cellin_2_5(2) <= cellout_1_5(2);cellin_2_4(0) <= cellout_1_4(0);cellin_2_4(1) <= cellout_1_4(1);cellin_2_4(2) <= cellout_1_4(2);cellin_2_4(3) <= cellout_1_4(3);cellin_2_3(0) <= cellout_1_3(0);cellin_2_3(1) <= cellout_1_3(1);cellin_2_3(2) <= cellout_1_3(2);cellin_2_3(3) <= cellout_1_3(3);cellin_2_2(0) <= cellout_1_2(0);cellin_2_2(1) <= cellout_1_2(1);cellin_2_2(2) <= cellout_1_2(2);cellin_2_2(3) <= cellout_1_2(3);cellin_2_1(0) <= cellout_1_1(0);cellin_2_1(1) <= cellout_1_1(1);cellin_2_1(2) <= cellout_1_1(2);cellin_2_1(3) <= cellout_1_1(3);cellin_4_10(0) <= cellout_3_10(0);cellin_4_9(0) <= cellout_3_9(0);cellin_4_9(1) <= cellout_3_9(1);cellin_4_8(0) <= cellout_3_8(0);cellin_4_7(0) <= cellout_3_7(0);cellin_4_6(0) <= cellout_3_6(0);cellin_4_5(0) <= cellout_3_5(0);cellin_4_5(1) <= cellout_3_5(1);cellin_4_4(0) <= cellout_3_4(0);cellin_4_4(1) <= cellout_3_4(1);cellin_4_3(0) <= cellout_3_3(0);cellin_4_3(1) <= cellout_3_3(1);cellin_4_2(0) <= cellout_3_2(0);cellin_4_2(1) <= cellout_3_2(1);cellin_4_1(0) <= cellout_3_1(0);cellin_4_1(1) <= cellout_3_1(1);cellin_6_11(0) <= cellout_5_11(0);cellin_6_10(0) <= cellout_5_10(0);cellin_6_10(1) <= cellout_5_10(1);cellin_6_9(0) <= cellout_5_9(0);cellin_6_9(1) <= cellout_5_9(1);cellin_6_8(0) <= cellout_5_8(0);cellin_6_8(1) <= cellout_5_8(1);cellin_6_7(0) <= cellout_5_7(0);cellin_6_7(1) <= cellout_5_7(1);cellin_6_6(0) <= cellout_5_6(0);cellin_6_6(1) <= cellout_5_6(1);cellin_6_5(0) <= cellout_5_5(0);cellin_6_5(1) <= cellout_5_5(1);cellin_6_4(0) <= cellout_5_4(0);cellin_6_4(1) <= cellout_5_4(1);cellin_6_3(0) <= cellout_5_3(0);cellin_6_3(1) <= cellout_5_3(1);cellin_6_3(2) <= cellout_5_3(2);cellin_6_2(0) <= cellout_5_2(0);cellin_6_2(1) <= cellout_5_2(1);cellin_6_1(0) <= cellout_5_1(0);cellin_6_1(1) <= cellout_5_1(1);cellin_8_11(0) <= cellout_7_11(0);cellin_8_10(0) <= cellout_7_10(0);cellin_8_10(1) <= cellout_7_10(1);cellin_8_9(0) <= cellout_7_9(0);cellin_8_9(1) <= cellout_7_9(1);cellin_8_8(0) <= cellout_7_8(0);cellin_8_7(0) <= cellout_7_7(0);cellin_8_7(1) <= cellout_7_7(1);cellin_8_6(0) <= cellout_7_6(0);cellin_8_6(1) <= cellout_7_6(1);cellin_8_5(0) <= cellout_7_5(0);cellin_8_5(1) <= cellout_7_5(1);cellin_8_4(0) <= cellout_7_4(0);cellin_8_4(1) <= cellout_7_4(1);cellin_8_3(0) <= cellout_7_3(0);cellin_8_3(1) <= cellout_7_3(1);cellin_8_2(0) <= cellout_7_2(0);cellin_8_2(1) <= cellout_7_2(1);cellin_8_1(0) <= cellout_7_1(0);cellin_8_1(1) <= cellout_7_1(1);cellin_10_11(0) <= cellout_9_11(0);cellin_10_11(1) <= cellout_9_11(1);cellin_10_10(0) <= cellout_9_10(0);cellin_10_9(0) <= cellout_9_9(0);cellin_10_9(1) <= cellout_9_9(1);cellin_10_9(2) <= cellout_9_9(2);cellin_10_8(0) <= cellout_9_8(0);cellin_10_8(1) <= cellout_9_8(1);cellin_10_7(0) <= cellout_9_7(0);cellin_10_7(1) <= cellout_9_7(1);cellin_10_7(2) <= cellout_9_7(2);cellin_10_6(0) <= cellout_9_6(0);cellin_10_6(1) <= cellout_9_6(1);cellin_10_6(2) <= cellout_9_6(2);cellin_10_5(0) <= cellout_9_5(0);cellin_10_5(1) <= cellout_9_5(1);cellin_10_4(0) <= cellout_9_4(0);cellin_10_4(1) <= cellout_9_4(1);cellin_10_3(0) <= cellout_9_3(0);cellin_10_3(1) <= cellout_9_3(1);cellin_10_3(2) <= cellout_9_3(2);cellin_10_2(0) <= cellout_9_2(0);cellin_10_2(1) <= cellout_9_2(1);cellin_10_1(0) <= cellout_9_1(0);cellin_10_1(1) <= cellout_9_1(1);cellin_12_11(0) <= cellout_11_11(0);cellin_12_11(1) <= cellout_11_11(1);cellin_12_10(0) <= cellout_11_10(0);cellin_12_9(0) <= cellout_11_9(0);cellin_12_8(0) <= cellout_11_8(0);cellin_12_8(1) <= cellout_11_8(1);cellin_12_7(0) <= cellout_11_7(0);cellin_12_7(1) <= cellout_11_7(1);cellin_12_6(0) <= cellout_11_6(0);cellin_12_6(1) <= cellout_11_6(1);cellin_12_5(0) <= cellout_11_5(0);cellin_12_5(1) <= cellout_11_5(1);cellin_12_4(0) <= cellout_11_4(0);cellin_12_4(1) <= cellout_11_4(1);cellin_12_3(0) <= cellout_11_3(0);cellin_12_3(1) <= cellout_11_3(1);cellin_12_2(0) <= cellout_11_2(0);cellin_12_2(1) <= cellout_11_2(1);cellin_12_1(0) <= cellout_11_1(0);cellin_12_1(1) <= cellout_11_1(1);cellin_14_11(0) <= cellout_13_11(0);cellin_14_10(0) <= cellout_13_10(0);cellin_14_10(1) <= cellout_13_10(1);cellin_14_10(2) <= cellout_13_10(2);cellin_14_9(0) <= cellout_13_9(0);cellin_14_8(0) <= cellout_13_8(0);cellin_14_8(1) <= cellout_13_8(1);cellin_14_8(2) <= cellout_13_8(2);cellin_14_8(3) <= cellout_13_8(3);cellin_14_7(0) <= cellout_13_7(0);cellin_14_7(1) <= cellout_13_7(1);cellin_14_7(2) <= cellout_13_7(2);cellin_14_6(0) <= cellout_13_6(0);cellin_14_6(1) <= cellout_13_6(1);cellin_14_6(2) <= cellout_13_6(2);cellin_14_6(3) <= cellout_13_6(3);cellin_14_6(4) <= cellout_13_6(4);cellin_14_5(0) <= cellout_13_5(0);cellin_14_5(1) <= cellout_13_5(1);cellin_14_5(2) <= cellout_13_5(2);cellin_14_5(3) <= cellout_13_5(3);cellin_14_5(4) <= cellout_13_5(4);cellin_14_4(0) <= cellout_13_4(0);cellin_14_4(1) <= cellout_13_4(1);cellin_14_4(2) <= cellout_13_4(2);cellin_14_4(3) <= cellout_13_4(3);cellin_14_4(4) <= cellout_13_4(4);cellin_14_4(5) <= cellout_13_4(5);cellin_14_3(0) <= cellout_13_3(0);cellin_14_3(1) <= cellout_13_3(1);cellin_14_3(2) <= cellout_13_3(2);cellin_14_3(3) <= cellout_13_3(3);cellin_14_3(4) <= cellout_13_3(4);cellin_14_3(5) <= cellout_13_3(5);cellin_14_2(0) <= cellout_13_2(0);cellin_14_2(1) <= cellout_13_2(1);cellin_14_2(2) <= cellout_13_2(2);cellin_14_2(3) <= cellout_13_2(3);cellin_14_2(4) <= cellout_13_2(4);cellin_14_2(5) <= cellout_13_2(5);cellin_14_1(0) <= cellout_13_1(0);cellin_14_1(1) <= cellout_13_1(1);cellin_14_1(2) <= cellout_13_1(2);cellin_14_1(3) <= cellout_13_1(3);cellin_14_1(4) <= cellout_13_1(4);cellin_14_1(5) <= cellout_13_1(5);cellin_16_11(0) <= cellout_15_11(0);cellin_16_10(0) <= cellout_15_10(0);cellin_16_9(0) <= cellout_15_9(0);cellin_16_8(0) <= cellout_15_8(0);cellin_16_8(1) <= cellout_15_8(1);cellin_16_8(2) <= cellout_15_8(2);cellin_16_7(0) <= cellout_15_7(0);cellin_16_7(1) <= cellout_15_7(1);cellin_16_6(0) <= cellout_15_6(0);cellin_16_6(1) <= cellout_15_6(1);cellin_16_5(0) <= cellout_15_5(0);cellin_16_5(1) <= cellout_15_5(1);cellin_16_5(2) <= cellout_15_5(2);cellin_16_4(0) <= cellout_15_4(0);cellin_16_4(1) <= cellout_15_4(1);cellin_16_3(0) <= cellout_15_3(0);cellin_16_3(1) <= cellout_15_3(1);cellin_16_3(2) <= cellout_15_3(2);cellin_16_2(0) <= cellout_15_2(0);cellin_16_2(1) <= cellout_15_2(1);cellin_16_2(2) <= cellout_15_2(2);cellin_16_1(0) <= cellout_15_1(0);cellin_16_1(1) <= cellout_15_1(1);cellin_16_1(2) <= cellout_15_1(2);out_1 <= cellin_17_1;out_2 <= cellin_17_2;out_3 <= cellin_17_3;out_4 <= cellin_17_4;out_5 <= cellin_17_5;out_6 <= cellin_17_6;out_7 <= cellin_17_7;out_8 <= cellin_17_8;out_9 <= cellin_17_9;out_10 <= cellin_17_10;out_11 <= cellin_17_11;end generated;