library ieee;use ieee.std_logic_1164.all;entity fir_cs isport (  clk, reset : in std_logic;  in_1_4 : in std_logic_vector(3 downto 0);  in_1_5 : in std_logic_vector(7 downto 0);  in_1_6 : in std_logic_vector(13 downto 0);  in_1_7 : in std_logic_vector(17 downto 0);  in_1_8 : in std_logic_vector(13 downto 0);  in_1_9 : in std_logic_vector(9 downto 0);  in_1_10 : in std_logic_vector(3 downto 0);  out_2 : out std_logic_vector(1 downto 0);  out_3 : out std_logic_vector(1 downto 0);  out_4 : out std_logic_vector(1 downto 0);  out_5 : out std_logic_vector(1 downto 0);  out_6 : out std_logic_vector(1 downto 0);  out_7 : out std_logic_vector(0 downto 0);  out_8 : out std_logic_vector(0 downto 0);  out_9 : out std_logic_vector(0 downto 0);  out_10 : out std_logic_vector(0 downto 0));end fir_cs;architecture generated of fir_cs iscomponent faport (in1, in2, in3 : in  std_logic;      outs, outc    : out std_logic);end component;component haport (in1, in2   : in  std_logic;      outs, outc : out std_logic);end component;component fa_nocport (in1, in2, in3 : in  std_logic;      outs          : out std_logic);end component;component ha_nocport (in1, in2 : in  std_logic;      outs     : out std_logic);end component;component dffport (clk, reset : in std_logic;      d : in  std_logic;      q : out std_logic);end component;signal cellin_1_4 : std_logic_vector(3 downto 0);signal cellin_1_5 : std_logic_vector(7 downto 0);signal cellin_1_6 : std_logic_vector(13 downto 0);signal cellin_1_7 : std_logic_vector(17 downto 0);signal cellin_1_8 : std_logic_vector(13 downto 0);signal cellin_1_9 : std_logic_vector(9 downto 0);signal cellin_1_10 : std_logic_vector(3 downto 0);signal cellin_2_3 : std_logic_vector(0 downto 0);signal cellin_2_4 : std_logic_vector(3 downto 0);signal cellin_2_5 : std_logic_vector(7 downto 0);signal cellin_2_6 : std_logic_vector(11 downto 0);signal cellin_2_7 : std_logic_vector(9 downto 0);signal cellin_2_8 : std_logic_vector(8 downto 0);signal cellin_2_9 : std_logic_vector(4 downto 0);signal cellin_2_10 : std_logic_vector(1 downto 0);signal cellin_3_3 : std_logic_vector(1 downto 0);signal cellin_3_4 : std_logic_vector(3 downto 0);signal cellin_3_5 : std_logic_vector(7 downto 0);signal cellin_3_6 : std_logic_vector(6 downto 0);signal cellin_3_7 : std_logic_vector(6 downto 0);signal cellin_3_8 : std_logic_vector(3 downto 0);signal cellin_3_9 : std_logic_vector(3 downto 0);signal cellin_3_10 : std_logic_vector(0 downto 0);signal cellin_4_3 : std_logic_vector(2 downto 0);signal cellin_4_4 : std_logic_vector(3 downto 0);signal cellin_4_5 : std_logic_vector(5 downto 0);signal cellin_4_6 : std_logic_vector(4 downto 0);signal cellin_4_7 : std_logic_vector(3 downto 0);signal cellin_4_8 : std_logic_vector(2 downto 0);signal cellin_4_9 : std_logic_vector(1 downto 0);signal cellin_4_10 : std_logic_vector(0 downto 0);signal cellin_5_2 : std_logic_vector(0 downto 0);signal cellin_5_3 : std_logic_vector(1 downto 0);signal cellin_5_4 : std_logic_vector(3 downto 0);signal cellin_5_5 : std_logic_vector(2 downto 0);signal cellin_5_6 : std_logic_vector(3 downto 0);signal cellin_5_7 : std_logic_vector(2 downto 0);signal cellin_5_8 : std_logic_vector(1 downto 0);signal cellin_5_9 : std_logic_vector(0 downto 0);signal cellin_5_10 : std_logic_vector(0 downto 0);signal cellin_6_2 : std_logic_vector(0 downto 0);signal cellin_6_3 : std_logic_vector(2 downto 0);signal cellin_6_4 : std_logic_vector(2 downto 0);signal cellin_6_5 : std_logic_vector(1 downto 0);signal cellin_6_6 : std_logic_vector(2 downto 0);signal cellin_6_7 : std_logic_vector(1 downto 0);signal cellin_6_8 : std_logic_vector(0 downto 0);signal cellin_6_9 : std_logic_vector(0 downto 0);signal cellin_6_10 : std_logic_vector(0 downto 0);signal cellin_7_2 : std_logic_vector(1 downto 0);signal cellin_7_3 : std_logic_vector(1 downto 0);signal cellin_7_4 : std_logic_vector(1 downto 0);signal cellin_7_5 : std_logic_vector(1 downto 0);signal cellin_7_6 : std_logic_vector(1 downto 0);signal cellin_7_7 : std_logic_vector(0 downto 0);signal cellin_7_8 : std_logic_vector(0 downto 0);signal cellin_7_9 : std_logic_vector(0 downto 0);signal cellin_7_10 : std_logic_vector(0 downto 0);signal cellout_1_3 : std_logic_vector(0 downto 0);signal cellout_1_4 : std_logic_vector(3 downto 0);signal cellout_1_5 : std_logic_vector(7 downto 0);signal cellout_1_6 : std_logic_vector(11 downto 0);signal cellout_1_7 : std_logic_vector(9 downto 0);signal cellout_1_8 : std_logic_vector(8 downto 0);signal cellout_1_9 : std_logic_vector(4 downto 0);signal cellout_1_10 : std_logic_vector(1 downto 0);signal cellout_2_3 : std_logic_vector(1 downto 0);signal cellout_2_4 : std_logic_vector(3 downto 0);signal cellout_2_5 : std_logic_vector(7 downto 0);signal cellout_2_6 : std_logic_vector(6 downto 0);signal cellout_2_7 : std_logic_vector(6 downto 0);signal cellout_2_8 : std_logic_vector(3 downto 0);signal cellout_2_9 : std_logic_vector(3 downto 0);signal cellout_2_10 : std_logic_vector(0 downto 0);signal cellout_3_3 : std_logic_vector(2 downto 0);signal cellout_3_4 : std_logic_vector(3 downto 0);signal cellout_3_5 : std_logic_vector(5 downto 0);signal cellout_3_6 : std_logic_vector(4 downto 0);signal cellout_3_7 : std_logic_vector(3 downto 0);signal cellout_3_8 : std_logic_vector(2 downto 0);signal cellout_3_9 : std_logic_vector(1 downto 0);signal cellout_3_10 : std_logic_vector(0 downto 0);signal cellout_4_2 : std_logic_vector(0 downto 0);signal cellout_4_3 : std_logic_vector(1 downto 0);signal cellout_4_4 : std_logic_vector(3 downto 0);signal cellout_4_5 : std_logic_vector(2 downto 0);signal cellout_4_6 : std_logic_vector(3 downto 0);signal cellout_4_7 : std_logic_vector(2 downto 0);signal cellout_4_8 : std_logic_vector(1 downto 0);signal cellout_4_9 : std_logic_vector(0 downto 0);signal cellout_4_10 : std_logic_vector(0 downto 0);signal cellout_5_2 : std_logic_vector(0 downto 0);signal cellout_5_3 : std_logic_vector(2 downto 0);signal cellout_5_4 : std_logic_vector(2 downto 0);signal cellout_5_5 : std_logic_vector(1 downto 0);signal cellout_5_6 : std_logic_vector(2 downto 0);signal cellout_5_7 : std_logic_vector(1 downto 0);signal cellout_5_8 : std_logic_vector(0 downto 0);signal cellout_5_9 : std_logic_vector(0 downto 0);signal cellout_5_10 : std_logic_vector(0 downto 0);signal cellout_6_2 : std_logic_vector(1 downto 0);signal cellout_6_3 : std_logic_vector(1 downto 0);signal cellout_6_4 : std_logic_vector(1 downto 0);signal cellout_6_5 : std_logic_vector(1 downto 0);signal cellout_6_6 : std_logic_vector(1 downto 0);signal cellout_6_7 : std_logic_vector(0 downto 0);signal cellout_6_8 : std_logic_vector(0 downto 0);signal cellout_6_9 : std_logic_vector(0 downto 0);signal cellout_6_10 : std_logic_vector(0 downto 0);begincellin_1_10(0) <= in_1_10(0);cellin_1_10(1) <= in_1_10(1);cellin_1_10(2) <= in_1_10(2);cellin_1_10(3) <= in_1_10(3);cellin_1_9(0) <= in_1_9(0);cellin_1_9(1) <= in_1_9(1);cellin_1_9(2) <= in_1_9(2);cellin_1_9(3) <= in_1_9(3);cellin_1_9(4) <= in_1_9(4);cellin_1_9(5) <= in_1_9(5);cellin_1_9(6) <= in_1_9(6);cellin_1_9(7) <= in_1_9(7);cellin_1_9(8) <= in_1_9(8);cellin_1_9(9) <= in_1_9(9);cellin_1_8(0) <= in_1_8(0);cellin_1_8(1) <= in_1_8(1);cellin_1_8(2) <= in_1_8(2);cellin_1_8(3) <= in_1_8(3);cellin_1_8(4) <= in_1_8(4);cellin_1_8(5) <= in_1_8(5);cellin_1_8(6) <= in_1_8(6);cellin_1_8(7) <= in_1_8(7);cellin_1_8(8) <= in_1_8(8);cellin_1_8(9) <= in_1_8(9);cellin_1_8(10) <= in_1_8(10);cellin_1_8(11) <= in_1_8(11);cellin_1_8(12) <= in_1_8(12);cellin_1_8(13) <= in_1_8(13);cellin_1_7(0) <= in_1_7(0);cellin_1_7(1) <= in_1_7(1);cellin_1_7(2) <= in_1_7(2);cellin_1_7(3) <= in_1_7(3);cellin_1_7(4) <= in_1_7(4);cellin_1_7(5) <= in_1_7(5);cellin_1_7(6) <= in_1_7(6);cellin_1_7(7) <= in_1_7(7);cellin_1_7(8) <= in_1_7(8);cellin_1_7(9) <= in_1_7(9);cellin_1_7(10) <= in_1_7(10);cellin_1_7(11) <= in_1_7(11);cellin_1_7(12) <= in_1_7(12);cellin_1_7(13) <= in_1_7(13);cellin_1_7(14) <= in_1_7(14);cellin_1_7(15) <= in_1_7(15);cellin_1_7(16) <= in_1_7(16);cellin_1_7(17) <= in_1_7(17);cellin_1_6(0) <= in_1_6(0);cellin_1_6(1) <= in_1_6(1);cellin_1_6(2) <= in_1_6(2);cellin_1_6(3) <= in_1_6(3);cellin_1_6(4) <= in_1_6(4);cellin_1_6(5) <= in_1_6(5);cellin_1_6(6) <= in_1_6(6);cellin_1_6(7) <= in_1_6(7);cellin_1_6(8) <= in_1_6(8);cellin_1_6(9) <= in_1_6(9);cellin_1_6(10) <= in_1_6(10);cellin_1_6(11) <= in_1_6(11);cellin_1_6(12) <= in_1_6(12);cellin_1_6(13) <= in_1_6(13);cellin_1_5(0) <= in_1_5(0);cellin_1_5(1) <= in_1_5(1);cellin_1_5(2) <= in_1_5(2);cellin_1_5(3) <= in_1_5(3);cellin_1_5(4) <= in_1_5(4);cellin_1_5(5) <= in_1_5(5);cellin_1_5(6) <= in_1_5(6);cellin_1_5(7) <= in_1_5(7);cellin_1_4(0) <= in_1_4(0);cellin_1_4(1) <= in_1_4(1);cellin_1_4(2) <= in_1_4(2);cellin_1_4(3) <= in_1_4(3);add_1_10_3_2_1: fa port map(cellin_1_10(3), cellin_1_10(2), cellin_1_10(1), cellout_1_10(0), cellout_1_9(0));add_1_9_9_8_7: fa port map(cellin_1_9(9), cellin_1_9(8), cellin_1_9(7), cellout_1_9(1), cellout_1_8(0));add_1_9_6_5_4: fa port map(cellin_1_9(6), cellin_1_9(5), cellin_1_9(4), cellout_1_9(2), cellout_1_8(1));add_1_9_3_2_1: fa port map(cellin_1_9(3), cellin_1_9(2), cellin_1_9(1), cellout_1_9(3), cellout_1_8(2));add_1_8_13_12_11: fa port map(cellin_1_8(13), cellin_1_8(12), cellin_1_8(11), cellout_1_8(3), cellout_1_7(0));add_1_8_10_9_8: fa port map(cellin_1_8(10), cellin_1_8(9), cellin_1_8(8), cellout_1_8(4), cellout_1_7(1));add_1_8_7_6_5: fa port map(cellin_1_8(7), cellin_1_8(6), cellin_1_8(5), cellout_1_8(5), cellout_1_7(2));add_1_8_4_3_2: fa port map(cellin_1_8(4), cellin_1_8(3), cellin_1_8(2), cellout_1_8(6), cellout_1_7(3));add_1_7_17_16_15: fa port map(cellin_1_7(17), cellin_1_7(16), cellin_1_7(15), cellout_1_7(4), cellout_1_6(0));add_1_7_14_13_12: fa port map(cellin_1_7(14), cellin_1_7(13), cellin_1_7(12), cellout_1_7(5), cellout_1_6(1));add_1_7_11_10_9: fa port map(cellin_1_7(11), cellin_1_7(10), cellin_1_7(9), cellout_1_7(6), cellout_1_6(2));add_1_7_8_7_6: fa port map(cellin_1_7(8), cellin_1_7(7), cellin_1_7(6), cellout_1_7(7), cellout_1_6(3));add_1_7_5_4_3: fa port map(cellin_1_7(5), cellin_1_7(4), cellin_1_7(3), cellout_1_7(8), cellout_1_6(4));add_1_7_2_1_0: fa port map(cellin_1_7(2), cellin_1_7(1), cellin_1_7(0), cellout_1_7(9), cellout_1_6(5));add_1_6_13_12_11: fa port map(cellin_1_6(13), cellin_1_6(12), cellin_1_6(11), cellout_1_6(6), cellout_1_5(0));add_1_6_10_9_8: fa port map(cellin_1_6(10), cellin_1_6(9), cellin_1_6(8), cellout_1_6(7), cellout_1_5(1));add_1_6_7_6_5: fa port map(cellin_1_6(7), cellin_1_6(6), cellin_1_6(5), cellout_1_6(8), cellout_1_5(2));add_1_6_4_3_2: fa port map(cellin_1_6(4), cellin_1_6(3), cellin_1_6(2), cellout_1_6(9), cellout_1_5(3));add_1_5_7_6_5: fa port map(cellin_1_5(7), cellin_1_5(6), cellin_1_5(5), cellout_1_5(4), cellout_1_4(0));add_1_5_4_3_2: fa port map(cellin_1_5(4), cellin_1_5(3), cellin_1_5(2), cellout_1_5(5), cellout_1_4(1));add_1_4_3_2_1: fa port map(cellin_1_4(3), cellin_1_4(2), cellin_1_4(1), cellout_1_4(2), cellout_1_3(0));add_2_9_4_3_2: fa port map(cellin_2_9(4), cellin_2_9(3), cellin_2_9(2), cellout_2_9(1), cellout_2_8(0));add_2_8_8_7_6: fa port map(cellin_2_8(8), cellin_2_8(7), cellin_2_8(6), cellout_2_8(1), cellout_2_7(0));add_2_8_5_4_3: fa port map(cellin_2_8(5), cellin_2_8(4), cellin_2_8(3), cellout_2_8(2), cellout_2_7(1));add_2_8_2_1_0: fa port map(cellin_2_8(2), cellin_2_8(1), cellin_2_8(0), cellout_2_8(3), cellout_2_7(2));add_2_7_9_8_7: fa port map(cellin_2_7(9), cellin_2_7(8), cellin_2_7(7), cellout_2_7(3), cellout_2_6(0));add_2_7_6_5_4: fa port map(cellin_2_7(6), cellin_2_7(5), cellin_2_7(4), cellout_2_7(4), cellout_2_6(1));add_2_7_3_2_1: fa port map(cellin_2_7(3), cellin_2_7(2), cellin_2_7(1), cellout_2_7(5), cellout_2_6(2));add_2_6_11_10_9: fa port map(cellin_2_6(11), cellin_2_6(10), cellin_2_6(9), cellout_2_6(3), cellout_2_5(0));add_2_6_8_7_6: fa port map(cellin_2_6(8), cellin_2_6(7), cellin_2_6(6), cellout_2_6(4), cellout_2_5(1));add_2_6_5_4_3: fa port map(cellin_2_6(5), cellin_2_6(4), cellin_2_6(3), cellout_2_6(5), cellout_2_5(2));add_2_6_2_1_0: fa port map(cellin_2_6(2), cellin_2_6(1), cellin_2_6(0), cellout_2_6(6), cellout_2_5(3));add_2_5_7_6_5: fa port map(cellin_2_5(7), cellin_2_5(6), cellin_2_5(5), cellout_2_5(4), cellout_2_4(0));add_2_5_4_3_2: fa port map(cellin_2_5(4), cellin_2_5(3), cellin_2_5(2), cellout_2_5(5), cellout_2_4(1));add_2_4_3_2_1: fa port map(cellin_2_4(3), cellin_2_4(2), cellin_2_4(1), cellout_2_4(2), cellout_2_3(0));add_3_9_3_2_1: fa port map(cellin_3_9(3), cellin_3_9(2), cellin_3_9(1), cellout_3_9(0), cellout_3_8(0));add_3_8_3_2_1: fa port map(cellin_3_8(3), cellin_3_8(2), cellin_3_8(1), cellout_3_8(1), cellout_3_7(0));add_3_7_6_5_4: fa port map(cellin_3_7(6), cellin_3_7(5), cellin_3_7(4), cellout_3_7(1), cellout_3_6(0));add_3_7_3_2_1: fa port map(cellin_3_7(3), cellin_3_7(2), cellin_3_7(1), cellout_3_7(2), cellout_3_6(1));add_3_6_6_5_4: fa port map(cellin_3_6(6), cellin_3_6(5), cellin_3_6(4), cellout_3_6(2), cellout_3_5(0));add_3_6_3_2_1: fa port map(cellin_3_6(3), cellin_3_6(2), cellin_3_6(1), cellout_3_6(3), cellout_3_5(1));add_3_5_7_6_5: fa port map(cellin_3_5(7), cellin_3_5(6), cellin_3_5(5), cellout_3_5(2), cellout_3_4(0));add_3_5_4_3_2: fa port map(cellin_3_5(4), cellin_3_5(3), cellin_3_5(2), cellout_3_5(3), cellout_3_4(1));add_3_4_3_2_1: fa port map(cellin_3_4(3), cellin_3_4(2), cellin_3_4(1), cellout_3_4(2), cellout_3_3(0));add_4_8_2_1_0: fa port map(cellin_4_8(2), cellin_4_8(1), cellin_4_8(0), cellout_4_8(1), cellout_4_7(0));add_4_7_3_2_1: fa port map(cellin_4_7(3), cellin_4_7(2), cellin_4_7(1), cellout_4_7(1), cellout_4_6(0));add_4_6_4_3_2: fa port map(cellin_4_6(4), cellin_4_6(3), cellin_4_6(2), cellout_4_6(1), cellout_4_5(0));add_4_5_5_4_3: fa port map(cellin_4_5(5), cellin_4_5(4), cellin_4_5(3), cellout_4_5(1), cellout_4_4(0));add_4_5_2_1_0: fa port map(cellin_4_5(2), cellin_4_5(1), cellin_4_5(0), cellout_4_5(2), cellout_4_4(1));add_4_4_3_2_1: fa port map(cellin_4_4(3), cellin_4_4(2), cellin_4_4(1), cellout_4_4(2), cellout_4_3(0));add_4_3_2_1_0: fa port map(cellin_4_3(2), cellin_4_3(1), cellin_4_3(0), cellout_4_3(1), cellout_4_2(0));add_5_7_2_1_0: fa port map(cellin_5_7(2), cellin_5_7(1), cellin_5_7(0), cellout_5_7(1), cellout_5_6(0));add_5_6_3_2_1: fa port map(cellin_5_6(3), cellin_5_6(2), cellin_5_6(1), cellout_5_6(1), cellout_5_5(0));add_5_5_2_1_0: fa port map(cellin_5_5(2), cellin_5_5(1), cellin_5_5(0), cellout_5_5(1), cellout_5_4(0));add_5_4_3_2_1: fa port map(cellin_5_4(3), cellin_5_4(2), cellin_5_4(1), cellout_5_4(1), cellout_5_3(0));add_6_6_2_1_0: fa port map(cellin_6_6(2), cellin_6_6(1), cellin_6_6(0), cellout_6_6(1), cellout_6_5(0));add_6_4_2_1_0: fa port map(cellin_6_4(2), cellin_6_4(1), cellin_6_4(0), cellout_6_4(1), cellout_6_3(0));add_6_3_2_1_0: fa port map(cellin_6_3(2), cellin_6_3(1), cellin_6_3(0), cellout_6_3(1), cellout_6_2(0));add_2_10_1_0: ha port map(cellin_2_10(1), cellin_2_10(0), cellout_2_10(0), cellout_2_9(0));add_4_9_1_0: ha port map(cellin_4_9(1), cellin_4_9(0), cellout_4_9(0), cellout_4_8(0));add_5_8_1_0: ha port map(cellin_5_8(1), cellin_5_8(0), cellout_5_8(0), cellout_5_7(0));add_6_7_1_0: ha port map(cellin_6_7(1), cellin_6_7(0), cellout_6_7(0), cellout_6_6(0));add_6_5_1_0: ha port map(cellin_6_5(1), cellin_6_5(0), cellout_6_5(1), cellout_6_4(0));cellout_1_10(1) <= cellin_1_10(0);cellout_1_9(4) <= cellin_1_9(0);cellout_1_8(7) <= cellin_1_8(1);cellout_1_8(8) <= cellin_1_8(0);cellout_1_6(10) <= cellin_1_6(1);cellout_1_6(11) <= cellin_1_6(0);cellout_1_5(6) <= cellin_1_5(1);cellout_1_5(7) <= cellin_1_5(0);cellout_1_4(3) <= cellin_1_4(0);cellout_2_9(2) <= cellin_2_9(1);cellout_2_9(3) <= cellin_2_9(0);cellout_2_7(6) <= cellin_2_7(0);cellout_2_5(6) <= cellin_2_5(1);cellout_2_5(7) <= cellin_2_5(0);cellout_2_4(3) <= cellin_2_4(0);cellout_2_3(1) <= cellin_2_3(0);cellout_3_10(0) <= cellin_3_10(0);cellout_3_9(1) <= cellin_3_9(0);cellout_3_8(2) <= cellin_3_8(0);cellout_3_7(3) <= cellin_3_7(0);cellout_3_6(4) <= cellin_3_6(0);cellout_3_5(4) <= cellin_3_5(1);cellout_3_5(5) <= cellin_3_5(0);cellout_3_4(3) <= cellin_3_4(0);cellout_3_3(1) <= cellin_3_3(1);cellout_3_3(2) <= cellin_3_3(0);cellout_4_10(0) <= cellin_4_10(0);cellout_4_7(2) <= cellin_4_7(0);cellout_4_6(2) <= cellin_4_6(1);cellout_4_6(3) <= cellin_4_6(0);cellout_4_4(3) <= cellin_4_4(0);cellout_5_10(0) <= cellin_5_10(0);cellout_5_9(0) <= cellin_5_9(0);cellout_5_6(2) <= cellin_5_6(0);cellout_5_4(2) <= cellin_5_4(0);cellout_5_3(1) <= cellin_5_3(1);cellout_5_3(2) <= cellin_5_3(0);cellout_5_2(0) <= cellin_5_2(0);cellout_6_10(0) <= cellin_6_10(0);cellout_6_9(0) <= cellin_6_9(0);cellout_6_8(0) <= cellin_6_8(0);cellout_6_2(1) <= cellin_6_2(0);reg_3_10_0: dff port map(clk, reset, cellout_3_10(0), cellin_4_10(0));reg_3_9_0: dff port map(clk, reset, cellout_3_9(0), cellin_4_9(0));reg_3_9_1: dff port map(clk, reset, cellout_3_9(1), cellin_4_9(1));reg_3_8_0: dff port map(clk, reset, cellout_3_8(0), cellin_4_8(0));reg_3_8_1: dff port map(clk, reset, cellout_3_8(1), cellin_4_8(1));reg_3_8_2: dff port map(clk, reset, cellout_3_8(2), cellin_4_8(2));reg_3_7_0: dff port map(clk, reset, cellout_3_7(0), cellin_4_7(0));reg_3_7_1: dff port map(clk, reset, cellout_3_7(1), cellin_4_7(1));reg_3_7_2: dff port map(clk, reset, cellout_3_7(2), cellin_4_7(2));reg_3_7_3: dff port map(clk, reset, cellout_3_7(3), cellin_4_7(3));reg_3_6_0: dff port map(clk, reset, cellout_3_6(0), cellin_4_6(0));reg_3_6_1: dff port map(clk, reset, cellout_3_6(1), cellin_4_6(1));reg_3_6_2: dff port map(clk, reset, cellout_3_6(2), cellin_4_6(2));reg_3_6_3: dff port map(clk, reset, cellout_3_6(3), cellin_4_6(3));reg_3_6_4: dff port map(clk, reset, cellout_3_6(4), cellin_4_6(4));reg_3_5_0: dff port map(clk, reset, cellout_3_5(0), cellin_4_5(0));reg_3_5_1: dff port map(clk, reset, cellout_3_5(1), cellin_4_5(1));reg_3_5_2: dff port map(clk, reset, cellout_3_5(2), cellin_4_5(2));reg_3_5_3: dff port map(clk, reset, cellout_3_5(3), cellin_4_5(3));reg_3_5_4: dff port map(clk, reset, cellout_3_5(4), cellin_4_5(4));reg_3_5_5: dff port map(clk, reset, cellout_3_5(5), cellin_4_5(5));reg_3_4_0: dff port map(clk, reset, cellout_3_4(0), cellin_4_4(0));reg_3_4_1: dff port map(clk, reset, cellout_3_4(1), cellin_4_4(1));reg_3_4_2: dff port map(clk, reset, cellout_3_4(2), cellin_4_4(2));reg_3_4_3: dff port map(clk, reset, cellout_3_4(3), cellin_4_4(3));reg_3_3_0: dff port map(clk, reset, cellout_3_3(0), cellin_4_3(0));reg_3_3_1: dff port map(clk, reset, cellout_3_3(1), cellin_4_3(1));reg_3_3_2: dff port map(clk, reset, cellout_3_3(2), cellin_4_3(2));reg_6_10_0: dff port map(clk, reset, cellout_6_10(0), cellin_7_10(0));reg_6_9_0: dff port map(clk, reset, cellout_6_9(0), cellin_7_9(0));reg_6_8_0: dff port map(clk, reset, cellout_6_8(0), cellin_7_8(0));reg_6_7_0: dff port map(clk, reset, cellout_6_7(0), cellin_7_7(0));reg_6_6_0: dff port map(clk, reset, cellout_6_6(0), cellin_7_6(0));reg_6_6_1: dff port map(clk, reset, cellout_6_6(1), cellin_7_6(1));reg_6_5_0: dff port map(clk, reset, cellout_6_5(0), cellin_7_5(0));reg_6_5_1: dff port map(clk, reset, cellout_6_5(1), cellin_7_5(1));reg_6_4_0: dff port map(clk, reset, cellout_6_4(0), cellin_7_4(0));reg_6_4_1: dff port map(clk, reset, cellout_6_4(1), cellin_7_4(1));reg_6_3_0: dff port map(clk, reset, cellout_6_3(0), cellin_7_3(0));reg_6_3_1: dff port map(clk, reset, cellout_6_3(1), cellin_7_3(1));reg_6_2_0: dff port map(clk, reset, cellout_6_2(0), cellin_7_2(0));reg_6_2_1: dff port map(clk, reset, cellout_6_2(1), cellin_7_2(1));cellin_2_10(0) <= cellout_1_10(0);cellin_2_10(1) <= cellout_1_10(1);cellin_2_9(0) <= cellout_1_9(0);cellin_2_9(1) <= cellout_1_9(1);cellin_2_9(2) <= cellout_1_9(2);cellin_2_9(3) <= cellout_1_9(3);cellin_2_9(4) <= cellout_1_9(4);cellin_2_8(0) <= cellout_1_8(0);cellin_2_8(1) <= cellout_1_8(1);cellin_2_8(2) <= cellout_1_8(2);cellin_2_8(3) <= cellout_1_8(3);cellin_2_8(4) <= cellout_1_8(4);cellin_2_8(5) <= cellout_1_8(5);cellin_2_8(6) <= cellout_1_8(6);cellin_2_8(7) <= cellout_1_8(7);cellin_2_8(8) <= cellout_1_8(8);cellin_2_7(0) <= cellout_1_7(0);cellin_2_7(1) <= cellout_1_7(1);cellin_2_7(2) <= cellout_1_7(2);cellin_2_7(3) <= cellout_1_7(3);cellin_2_7(4) <= cellout_1_7(4);cellin_2_7(5) <= cellout_1_7(5);cellin_2_7(6) <= cellout_1_7(6);cellin_2_7(7) <= cellout_1_7(7);cellin_2_7(8) <= cellout_1_7(8);cellin_2_7(9) <= cellout_1_7(9);cellin_2_6(0) <= cellout_1_6(0);cellin_2_6(1) <= cellout_1_6(1);cellin_2_6(2) <= cellout_1_6(2);cellin_2_6(3) <= cellout_1_6(3);cellin_2_6(4) <= cellout_1_6(4);cellin_2_6(5) <= cellout_1_6(5);cellin_2_6(6) <= cellout_1_6(6);cellin_2_6(7) <= cellout_1_6(7);cellin_2_6(8) <= cellout_1_6(8);cellin_2_6(9) <= cellout_1_6(9);cellin_2_6(10) <= cellout_1_6(10);cellin_2_6(11) <= cellout_1_6(11);cellin_2_5(0) <= cellout_1_5(0);cellin_2_5(1) <= cellout_1_5(1);cellin_2_5(2) <= cellout_1_5(2);cellin_2_5(3) <= cellout_1_5(3);cellin_2_5(4) <= cellout_1_5(4);cellin_2_5(5) <= cellout_1_5(5);cellin_2_5(6) <= cellout_1_5(6);cellin_2_5(7) <= cellout_1_5(7);cellin_2_4(0) <= cellout_1_4(0);cellin_2_4(1) <= cellout_1_4(1);cellin_2_4(2) <= cellout_1_4(2);cellin_2_4(3) <= cellout_1_4(3);cellin_2_3(0) <= cellout_1_3(0);cellin_3_10(0) <= cellout_2_10(0);cellin_3_9(0) <= cellout_2_9(0);cellin_3_9(1) <= cellout_2_9(1);cellin_3_9(2) <= cellout_2_9(2);cellin_3_9(3) <= cellout_2_9(3);cellin_3_8(0) <= cellout_2_8(0);cellin_3_8(1) <= cellout_2_8(1);cellin_3_8(2) <= cellout_2_8(2);cellin_3_8(3) <= cellout_2_8(3);cellin_3_7(0) <= cellout_2_7(0);cellin_3_7(1) <= cellout_2_7(1);cellin_3_7(2) <= cellout_2_7(2);cellin_3_7(3) <= cellout_2_7(3);cellin_3_7(4) <= cellout_2_7(4);cellin_3_7(5) <= cellout_2_7(5);cellin_3_7(6) <= cellout_2_7(6);cellin_3_6(0) <= cellout_2_6(0);cellin_3_6(1) <= cellout_2_6(1);cellin_3_6(2) <= cellout_2_6(2);cellin_3_6(3) <= cellout_2_6(3);cellin_3_6(4) <= cellout_2_6(4);cellin_3_6(5) <= cellout_2_6(5);cellin_3_6(6) <= cellout_2_6(6);cellin_3_5(0) <= cellout_2_5(0);cellin_3_5(1) <= cellout_2_5(1);cellin_3_5(2) <= cellout_2_5(2);cellin_3_5(3) <= cellout_2_5(3);cellin_3_5(4) <= cellout_2_5(4);cellin_3_5(5) <= cellout_2_5(5);cellin_3_5(6) <= cellout_2_5(6);cellin_3_5(7) <= cellout_2_5(7);cellin_3_4(0) <= cellout_2_4(0);cellin_3_4(1) <= cellout_2_4(1);cellin_3_4(2) <= cellout_2_4(2);cellin_3_4(3) <= cellout_2_4(3);cellin_3_3(0) <= cellout_2_3(0);cellin_3_3(1) <= cellout_2_3(1);cellin_5_10(0) <= cellout_4_10(0);cellin_5_9(0) <= cellout_4_9(0);cellin_5_8(0) <= cellout_4_8(0);cellin_5_8(1) <= cellout_4_8(1);cellin_5_7(0) <= cellout_4_7(0);cellin_5_7(1) <= cellout_4_7(1);cellin_5_7(2) <= cellout_4_7(2);cellin_5_6(0) <= cellout_4_6(0);cellin_5_6(1) <= cellout_4_6(1);cellin_5_6(2) <= cellout_4_6(2);cellin_5_6(3) <= cellout_4_6(3);cellin_5_5(0) <= cellout_4_5(0);cellin_5_5(1) <= cellout_4_5(1);cellin_5_5(2) <= cellout_4_5(2);cellin_5_4(0) <= cellout_4_4(0);cellin_5_4(1) <= cellout_4_4(1);cellin_5_4(2) <= cellout_4_4(2);cellin_5_4(3) <= cellout_4_4(3);cellin_5_3(0) <= cellout_4_3(0);cellin_5_3(1) <= cellout_4_3(1);cellin_5_2(0) <= cellout_4_2(0);cellin_6_10(0) <= cellout_5_10(0);cellin_6_9(0) <= cellout_5_9(0);cellin_6_8(0) <= cellout_5_8(0);cellin_6_7(0) <= cellout_5_7(0);cellin_6_7(1) <= cellout_5_7(1);cellin_6_6(0) <= cellout_5_6(0);cellin_6_6(1) <= cellout_5_6(1);cellin_6_6(2) <= cellout_5_6(2);cellin_6_5(0) <= cellout_5_5(0);cellin_6_5(1) <= cellout_5_5(1);cellin_6_4(0) <= cellout_5_4(0);cellin_6_4(1) <= cellout_5_4(1);cellin_6_4(2) <= cellout_5_4(2);cellin_6_3(0) <= cellout_5_3(0);cellin_6_3(1) <= cellout_5_3(1);cellin_6_3(2) <= cellout_5_3(2);cellin_6_2(0) <= cellout_5_2(0);out_2 <= cellin_7_2;out_3 <= cellin_7_3;out_4 <= cellin_7_4;out_5 <= cellin_7_5;out_6 <= cellin_7_6;out_7 <= cellin_7_7;out_8 <= cellin_7_8;out_9 <= cellin_7_9;out_10 <= cellin_7_10;end generated;