library ieee;use ieee.std_logic_1164.all;entity fir_pp isport (clk, reset : in std_logic;  in_0 : in std_logic_vector(5 downto 0);  out_1_1 : out std_logic_vector(5 downto 0);  out_1_2 : out std_logic_vector(5 downto 0);  out_1_3 : out std_logic_vector(5 downto 0);  out_1_4 : out std_logic_vector(5 downto 0);  out_1_5 : out std_logic_vector(5 downto 0);  out_1_6 : out std_logic_vector(4 downto 0);  out_1_7 : out std_logic_vector(3 downto 0);  out_1_8 : out std_logic_vector(2 downto 0);  out_1_9 : out std_logic_vector(1 downto 0);  out_1_10 : out std_logic_vector(0 downto 0);  out_5_4 : out std_logic_vector(0 downto 0);  out_5_5 : out std_logic_vector(0 downto 0);  out_5_6 : out std_logic_vector(1 downto 0);  out_5_7 : out std_logic_vector(1 downto 0);  out_5_8 : out std_logic_vector(1 downto 0);  out_5_9 : out std_logic_vector(1 downto 0);  out_5_10 : out std_logic_vector(0 downto 0);  out_5_11 : out std_logic_vector(0 downto 0);  out_7_3 : out std_logic_vector(0 downto 0);  out_7_4 : out std_logic_vector(0 downto 0);  out_7_5 : out std_logic_vector(0 downto 0);  out_7_6 : out std_logic_vector(0 downto 0);  out_7_7 : out std_logic_vector(0 downto 0);  out_7_8 : out std_logic_vector(0 downto 0);  out_9_4 : out std_logic_vector(0 downto 0);  out_9_5 : out std_logic_vector(0 downto 0);  out_9_6 : out std_logic_vector(1 downto 0);  out_9_7 : out std_logic_vector(1 downto 0);  out_9_8 : out std_logic_vector(1 downto 0);  out_9_9 : out std_logic_vector(1 downto 0);  out_9_10 : out std_logic_vector(0 downto 0);  out_9_11 : out std_logic_vector(0 downto 0);  out_13_1 : out std_logic_vector(5 downto 0);  out_13_2 : out std_logic_vector(5 downto 0);  out_13_3 : out std_logic_vector(5 downto 0);  out_13_4 : out std_logic_vector(5 downto 0);  out_13_5 : out std_logic_vector(5 downto 0);  out_13_6 : out std_logic_vector(4 downto 0);  out_13_7 : out std_logic_vector(3 downto 0);  out_13_8 : out std_logic_vector(2 downto 0);  out_13_9 : out std_logic_vector(1 downto 0);  out_13_10 : out std_logic_vector(0 downto 0));end fir_pp;architecture generated of fir_pp isbeginout_1_1(0) <= in_0(0);out_1_1(1) <= in_0(1);out_1_1(2) <= in_0(2);out_1_1(3) <= in_0(3);out_1_1(4) <= in_0(4);out_1_1(5) <= not in_0(5);out_1_2(0) <= in_0(0);out_1_2(1) <= in_0(1);out_1_2(2) <= in_0(2);out_1_2(3) <= in_0(3);out_1_2(4) <= in_0(4);out_1_2(5) <= not in_0(5);out_1_3(0) <= in_0(0);out_1_3(1) <= in_0(1);out_1_3(2) <= in_0(2);out_1_3(3) <= in_0(3);out_1_3(4) <= in_0(4);out_1_3(5) <= not in_0(5);out_1_4(0) <= in_0(0);out_1_4(1) <= in_0(1);out_1_4(2) <= in_0(2);out_1_4(3) <= in_0(3);out_1_4(4) <= in_0(4);out_1_4(5) <= not in_0(5);out_1_5(0) <= in_0(0);out_1_5(1) <= in_0(1);out_1_5(2) <= in_0(2);out_1_5(3) <= in_0(3);out_1_5(4) <= in_0(4);out_1_5(5) <= not in_0(5);out_1_6(0) <= in_0(0);out_1_6(1) <= in_0(1);out_1_6(2) <= in_0(2);out_1_6(3) <= in_0(3);out_1_6(4) <= in_0(4);out_1_7(0) <= in_0(0);out_1_7(1) <= in_0(1);out_1_7(2) <= in_0(2);out_1_7(3) <= in_0(3);out_1_8(0) <= in_0(0);out_1_8(1) <= in_0(1);out_1_8(2) <= in_0(2);out_1_9(0) <= in_0(0);out_1_9(1) <= in_0(1);out_1_10(0) <= in_0(0);out_5_4(0) <= not in_0(5);out_5_5(0) <= in_0(4);out_5_6(0) <= in_0(3);out_5_6(1) <= not in_0(5);out_5_7(0) <= in_0(2);out_5_7(1) <= in_0(4);out_5_8(0) <= in_0(1);out_5_8(1) <= in_0(3);out_5_9(0) <= in_0(0);out_5_9(1) <= in_0(2);out_5_10(0) <= in_0(1);out_5_11(0) <= in_0(0);out_7_3(0) <= not in_0(5);out_7_4(0) <= in_0(4);out_7_5(0) <= in_0(3);out_7_6(0) <= in_0(2);out_7_7(0) <= in_0(1);out_7_8(0) <= in_0(0);out_9_4(0) <= not in_0(5);out_9_5(0) <= in_0(4);out_9_6(0) <= in_0(3);out_9_6(1) <= not in_0(5);out_9_7(0) <= in_0(2);out_9_7(1) <= in_0(4);out_9_8(0) <= in_0(1);out_9_8(1) <= in_0(3);out_9_9(0) <= in_0(0);out_9_9(1) <= in_0(2);out_9_10(0) <= in_0(1);out_9_11(0) <= in_0(0);out_13_1(0) <= in_0(0);out_13_1(1) <= in_0(1);out_13_1(2) <= in_0(2);out_13_1(3) <= in_0(3);out_13_1(4) <= in_0(4);out_13_1(5) <= not in_0(5);out_13_2(0) <= in_0(0);out_13_2(1) <= in_0(1);out_13_2(2) <= in_0(2);out_13_2(3) <= in_0(3);out_13_2(4) <= in_0(4);out_13_2(5) <= not in_0(5);out_13_3(0) <= in_0(0);out_13_3(1) <= in_0(1);out_13_3(2) <= in_0(2);out_13_3(3) <= in_0(3);out_13_3(4) <= in_0(4);out_13_3(5) <= not in_0(5);out_13_4(0) <= in_0(0);out_13_4(1) <= in_0(1);out_13_4(2) <= in_0(2);out_13_4(3) <= in_0(3);out_13_4(4) <= in_0(4);out_13_4(5) <= not in_0(5);out_13_5(0) <= in_0(0);out_13_5(1) <= in_0(1);out_13_5(2) <= in_0(2);out_13_5(3) <= in_0(3);out_13_5(4) <= in_0(4);out_13_5(5) <= not in_0(5);out_13_6(0) <= in_0(0);out_13_6(1) <= in_0(1);out_13_6(2) <= in_0(2);out_13_6(3) <= in_0(3);out_13_6(4) <= in_0(4);out_13_7(0) <= in_0(0);out_13_7(1) <= in_0(1);out_13_7(2) <= in_0(2);out_13_7(3) <= in_0(3);out_13_8(0) <= in_0(0);out_13_8(1) <= in_0(1);out_13_8(2) <= in_0(2);out_13_9(0) <= in_0(0);out_13_9(1) <= in_0(1);out_13_10(0) <= in_0(0);end generated;