library ieee;use ieee.std_logic_1164.all;entity fir_vma isport (  clk, reset : in std_logic;  in_1_2 : in std_logic_vector(1 downto 0);  in_1_3 : in std_logic_vector(1 downto 0);  in_1_4 : in std_logic_vector(1 downto 0);  in_1_5 : in std_logic_vector(1 downto 0);  in_1_6 : in std_logic_vector(1 downto 0);  in_1_7 : in std_logic_vector(0 downto 0);  in_1_8 : in std_logic_vector(0 downto 0);  in_1_9 : in std_logic_vector(0 downto 0);  in_1_10 : in std_logic_vector(0 downto 0);  out_1 : out std_logic_vector(0 downto 0);  out_2 : out std_logic_vector(0 downto 0);  out_3 : out std_logic_vector(0 downto 0);  out_4 : out std_logic_vector(0 downto 0);  out_5 : out std_logic_vector(0 downto 0);  out_6 : out std_logic_vector(0 downto 0);  out_7 : out std_logic_vector(0 downto 0);  out_8 : out std_logic_vector(0 downto 0);  out_9 : out std_logic_vector(0 downto 0);  out_10 : out std_logic_vector(0 downto 0));end fir_vma;architecture generated of fir_vma iscomponent faport (in1, in2, in3 : in  std_logic;      outs, outc    : out std_logic);end component;component haport (in1, in2   : in  std_logic;      outs, outc : out std_logic);end component;component fa_nocport (in1, in2, in3 : in  std_logic;      outs          : out std_logic);end component;component ha_nocport (in1, in2 : in  std_logic;      outs     : out std_logic);end component;component dffport (clk, reset : in std_logic;      d : in  std_logic;      q : out std_logic);end component;signal cellin_1_2 : std_logic_vector(1 downto 0);signal cellin_1_3 : std_logic_vector(1 downto 0);signal cellin_1_4 : std_logic_vector(1 downto 0);signal cellin_1_5 : std_logic_vector(1 downto 0);signal cellin_1_6 : std_logic_vector(1 downto 0);signal cellin_1_7 : std_logic_vector(0 downto 0);signal cellin_1_8 : std_logic_vector(0 downto 0);signal cellin_1_9 : std_logic_vector(0 downto 0);signal cellin_1_10 : std_logic_vector(0 downto 0);signal cellin_2_2 : std_logic_vector(1 downto 0);signal cellin_2_3 : std_logic_vector(1 downto 0);signal cellin_2_4 : std_logic_vector(1 downto 0);signal cellin_2_5 : std_logic_vector(2 downto 0);signal cellin_2_6 : std_logic_vector(0 downto 0);signal cellin_2_7 : std_logic_vector(0 downto 0);signal cellin_2_8 : std_logic_vector(0 downto 0);signal cellin_2_9 : std_logic_vector(0 downto 0);signal cellin_2_10 : std_logic_vector(0 downto 0);signal cellin_3_2 : std_logic_vector(1 downto 0);signal cellin_3_3 : std_logic_vector(1 downto 0);signal cellin_3_4 : std_logic_vector(2 downto 0);signal cellin_3_5 : std_logic_vector(0 downto 0);signal cellin_3_6 : std_logic_vector(0 downto 0);signal cellin_3_7 : std_logic_vector(0 downto 0);signal cellin_3_8 : std_logic_vector(0 downto 0);signal cellin_3_9 : std_logic_vector(0 downto 0);signal cellin_3_10 : std_logic_vector(0 downto 0);signal cellin_4_2 : std_logic_vector(1 downto 0);signal cellin_4_3 : std_logic_vector(2 downto 0);signal cellin_4_4 : std_logic_vector(0 downto 0);signal cellin_4_5 : std_logic_vector(0 downto 0);signal cellin_4_6 : std_logic_vector(0 downto 0);signal cellin_4_7 : std_logic_vector(0 downto 0);signal cellin_4_8 : std_logic_vector(0 downto 0);signal cellin_4_9 : std_logic_vector(0 downto 0);signal cellin_4_10 : std_logic_vector(0 downto 0);signal cellin_5_2 : std_logic_vector(2 downto 0);signal cellin_5_3 : std_logic_vector(0 downto 0);signal cellin_5_4 : std_logic_vector(0 downto 0);signal cellin_5_5 : std_logic_vector(0 downto 0);signal cellin_5_6 : std_logic_vector(0 downto 0);signal cellin_5_7 : std_logic_vector(0 downto 0);signal cellin_5_8 : std_logic_vector(0 downto 0);signal cellin_5_9 : std_logic_vector(0 downto 0);signal cellin_5_10 : std_logic_vector(0 downto 0);signal cellin_6_1 : std_logic_vector(0 downto 0);signal cellin_6_2 : std_logic_vector(0 downto 0);signal cellin_6_3 : std_logic_vector(0 downto 0);signal cellin_6_4 : std_logic_vector(0 downto 0);signal cellin_6_5 : std_logic_vector(0 downto 0);signal cellin_6_6 : std_logic_vector(0 downto 0);signal cellin_6_7 : std_logic_vector(0 downto 0);signal cellin_6_8 : std_logic_vector(0 downto 0);signal cellin_6_9 : std_logic_vector(0 downto 0);signal cellin_6_10 : std_logic_vector(0 downto 0);signal cellin_7_1 : std_logic_vector(0 downto 0);signal cellin_7_2 : std_logic_vector(0 downto 0);signal cellin_7_3 : std_logic_vector(0 downto 0);signal cellin_7_4 : std_logic_vector(0 downto 0);signal cellin_7_5 : std_logic_vector(0 downto 0);signal cellin_7_6 : std_logic_vector(0 downto 0);signal cellin_7_7 : std_logic_vector(0 downto 0);signal cellin_7_8 : std_logic_vector(0 downto 0);signal cellin_7_9 : std_logic_vector(0 downto 0);signal cellin_7_10 : std_logic_vector(0 downto 0);signal cellout_1_2 : std_logic_vector(1 downto 0);signal cellout_1_3 : std_logic_vector(1 downto 0);signal cellout_1_4 : std_logic_vector(1 downto 0);signal cellout_1_5 : std_logic_vector(2 downto 0);signal cellout_1_6 : std_logic_vector(0 downto 0);signal cellout_1_7 : std_logic_vector(0 downto 0);signal cellout_1_8 : std_logic_vector(0 downto 0);signal cellout_1_9 : std_logic_vector(0 downto 0);signal cellout_1_10 : std_logic_vector(0 downto 0);signal cellout_2_2 : std_logic_vector(1 downto 0);signal cellout_2_3 : std_logic_vector(1 downto 0);signal cellout_2_4 : std_logic_vector(2 downto 0);signal cellout_2_5 : std_logic_vector(0 downto 0);signal cellout_2_6 : std_logic_vector(0 downto 0);signal cellout_2_7 : std_logic_vector(0 downto 0);signal cellout_2_8 : std_logic_vector(0 downto 0);signal cellout_2_9 : std_logic_vector(0 downto 0);signal cellout_2_10 : std_logic_vector(0 downto 0);signal cellout_3_2 : std_logic_vector(1 downto 0);signal cellout_3_3 : std_logic_vector(2 downto 0);signal cellout_3_4 : std_logic_vector(0 downto 0);signal cellout_3_5 : std_logic_vector(0 downto 0);signal cellout_3_6 : std_logic_vector(0 downto 0);signal cellout_3_7 : std_logic_vector(0 downto 0);signal cellout_3_8 : std_logic_vector(0 downto 0);signal cellout_3_9 : std_logic_vector(0 downto 0);signal cellout_3_10 : std_logic_vector(0 downto 0);signal cellout_4_2 : std_logic_vector(2 downto 0);signal cellout_4_3 : std_logic_vector(0 downto 0);signal cellout_4_4 : std_logic_vector(0 downto 0);signal cellout_4_5 : std_logic_vector(0 downto 0);signal cellout_4_6 : std_logic_vector(0 downto 0);signal cellout_4_7 : std_logic_vector(0 downto 0);signal cellout_4_8 : std_logic_vector(0 downto 0);signal cellout_4_9 : std_logic_vector(0 downto 0);signal cellout_4_10 : std_logic_vector(0 downto 0);signal cellout_5_1 : std_logic_vector(0 downto 0);signal cellout_5_2 : std_logic_vector(0 downto 0);signal cellout_5_3 : std_logic_vector(0 downto 0);signal cellout_5_4 : std_logic_vector(0 downto 0);signal cellout_5_5 : std_logic_vector(0 downto 0);signal cellout_5_6 : std_logic_vector(0 downto 0);signal cellout_5_7 : std_logic_vector(0 downto 0);signal cellout_5_8 : std_logic_vector(0 downto 0);signal cellout_5_9 : std_logic_vector(0 downto 0);signal cellout_5_10 : std_logic_vector(0 downto 0);signal cellout_6_1 : std_logic_vector(0 downto 0);signal cellout_6_2 : std_logic_vector(0 downto 0);signal cellout_6_3 : std_logic_vector(0 downto 0);signal cellout_6_4 : std_logic_vector(0 downto 0);signal cellout_6_5 : std_logic_vector(0 downto 0);signal cellout_6_6 : std_logic_vector(0 downto 0);signal cellout_6_7 : std_logic_vector(0 downto 0);signal cellout_6_8 : std_logic_vector(0 downto 0);signal cellout_6_9 : std_logic_vector(0 downto 0);signal cellout_6_10 : std_logic_vector(0 downto 0);begincellin_1_10(0) <= in_1_10(0);cellin_1_9(0) <= in_1_9(0);cellin_1_8(0) <= in_1_8(0);cellin_1_7(0) <= in_1_7(0);cellin_1_6(0) <= in_1_6(0);cellin_1_6(1) <= in_1_6(1);cellin_1_5(0) <= in_1_5(0);cellin_1_5(1) <= in_1_5(1);cellin_1_4(0) <= in_1_4(0);cellin_1_4(1) <= in_1_4(1);cellin_1_3(0) <= in_1_3(0);cellin_1_3(1) <= in_1_3(1);cellin_1_2(0) <= in_1_2(0);cellin_1_2(1) <= in_1_2(1);add_2_5_2_1_0: fa port map(cellin_2_5(2), cellin_2_5(1), cellin_2_5(0), cellout_2_5(0), cellout_2_4(0));add_3_4_2_1_0: fa port map(cellin_3_4(2), cellin_3_4(1), cellin_3_4(0), cellout_3_4(0), cellout_3_3(0));add_4_3_2_1_0: fa port map(cellin_4_3(2), cellin_4_3(1), cellin_4_3(0), cellout_4_3(0), cellout_4_2(0));add_5_2_2_1_0: fa port map(cellin_5_2(2), cellin_5_2(1), cellin_5_2(0), cellout_5_2(0), cellout_5_1(0));add_1_6_1_0: ha port map(cellin_1_6(1), cellin_1_6(0), cellout_1_6(0), cellout_1_5(0));cellout_1_10(0) <= cellin_1_10(0);cellout_1_9(0) <= cellin_1_9(0);cellout_1_8(0) <= cellin_1_8(0);cellout_1_7(0) <= cellin_1_7(0);cellout_1_5(1) <= cellin_1_5(1);cellout_1_5(2) <= cellin_1_5(0);cellout_1_4(0) <= cellin_1_4(1);cellout_1_4(1) <= cellin_1_4(0);cellout_1_3(0) <= cellin_1_3(1);cellout_1_3(1) <= cellin_1_3(0);cellout_1_2(0) <= cellin_1_2(1);cellout_1_2(1) <= cellin_1_2(0);cellout_2_10(0) <= cellin_2_10(0);cellout_2_9(0) <= cellin_2_9(0);cellout_2_8(0) <= cellin_2_8(0);cellout_2_7(0) <= cellin_2_7(0);cellout_2_6(0) <= cellin_2_6(0);cellout_2_4(1) <= cellin_2_4(1);cellout_2_4(2) <= cellin_2_4(0);cellout_2_3(0) <= cellin_2_3(1);cellout_2_3(1) <= cellin_2_3(0);cellout_2_2(0) <= cellin_2_2(1);cellout_2_2(1) <= cellin_2_2(0);cellout_3_10(0) <= cellin_3_10(0);cellout_3_9(0) <= cellin_3_9(0);cellout_3_8(0) <= cellin_3_8(0);cellout_3_7(0) <= cellin_3_7(0);cellout_3_6(0) <= cellin_3_6(0);cellout_3_5(0) <= cellin_3_5(0);cellout_3_3(1) <= cellin_3_3(1);cellout_3_3(2) <= cellin_3_3(0);cellout_3_2(0) <= cellin_3_2(1);cellout_3_2(1) <= cellin_3_2(0);cellout_4_10(0) <= cellin_4_10(0);cellout_4_9(0) <= cellin_4_9(0);cellout_4_8(0) <= cellin_4_8(0);cellout_4_7(0) <= cellin_4_7(0);cellout_4_6(0) <= cellin_4_6(0);cellout_4_5(0) <= cellin_4_5(0);cellout_4_4(0) <= cellin_4_4(0);cellout_4_2(1) <= cellin_4_2(1);cellout_4_2(2) <= cellin_4_2(0);cellout_5_10(0) <= cellin_5_10(0);cellout_5_9(0) <= cellin_5_9(0);cellout_5_8(0) <= cellin_5_8(0);cellout_5_7(0) <= cellin_5_7(0);cellout_5_6(0) <= cellin_5_6(0);cellout_5_5(0) <= cellin_5_5(0);cellout_5_4(0) <= cellin_5_4(0);cellout_5_3(0) <= cellin_5_3(0);cellout_6_10(0) <= cellin_6_10(0);cellout_6_9(0) <= cellin_6_9(0);cellout_6_8(0) <= cellin_6_8(0);cellout_6_7(0) <= cellin_6_7(0);cellout_6_6(0) <= cellin_6_6(0);cellout_6_5(0) <= cellin_6_5(0);cellout_6_4(0) <= cellin_6_4(0);cellout_6_3(0) <= cellin_6_3(0);cellout_6_2(0) <= cellin_6_2(0);cellout_6_1(0) <= cellin_6_1(0);reg_3_10_0: dff port map(clk, reset, cellout_3_10(0), cellin_4_10(0));reg_3_9_0: dff port map(clk, reset, cellout_3_9(0), cellin_4_9(0));reg_3_8_0: dff port map(clk, reset, cellout_3_8(0), cellin_4_8(0));reg_3_7_0: dff port map(clk, reset, cellout_3_7(0), cellin_4_7(0));reg_3_6_0: dff port map(clk, reset, cellout_3_6(0), cellin_4_6(0));reg_3_5_0: dff port map(clk, reset, cellout_3_5(0), cellin_4_5(0));reg_3_4_0: dff port map(clk, reset, cellout_3_4(0), cellin_4_4(0));reg_3_3_0: dff port map(clk, reset, cellout_3_3(0), cellin_4_3(0));reg_3_3_1: dff port map(clk, reset, cellout_3_3(1), cellin_4_3(1));reg_3_3_2: dff port map(clk, reset, cellout_3_3(2), cellin_4_3(2));reg_3_2_0: dff port map(clk, reset, cellout_3_2(0), cellin_4_2(0));reg_3_2_1: dff port map(clk, reset, cellout_3_2(1), cellin_4_2(1));reg_6_10_0: dff port map(clk, reset, cellout_6_10(0), cellin_7_10(0));reg_6_9_0: dff port map(clk, reset, cellout_6_9(0), cellin_7_9(0));reg_6_8_0: dff port map(clk, reset, cellout_6_8(0), cellin_7_8(0));reg_6_7_0: dff port map(clk, reset, cellout_6_7(0), cellin_7_7(0));reg_6_6_0: dff port map(clk, reset, cellout_6_6(0), cellin_7_6(0));reg_6_5_0: dff port map(clk, reset, cellout_6_5(0), cellin_7_5(0));reg_6_4_0: dff port map(clk, reset, cellout_6_4(0), cellin_7_4(0));reg_6_3_0: dff port map(clk, reset, cellout_6_3(0), cellin_7_3(0));reg_6_2_0: dff port map(clk, reset, cellout_6_2(0), cellin_7_2(0));reg_6_1_0: dff port map(clk, reset, cellout_6_1(0), cellin_7_1(0));cellin_2_10(0) <= cellout_1_10(0);cellin_2_9(0) <= cellout_1_9(0);cellin_2_8(0) <= cellout_1_8(0);cellin_2_7(0) <= cellout_1_7(0);cellin_2_6(0) <= cellout_1_6(0);cellin_2_5(0) <= cellout_1_5(0);cellin_2_5(1) <= cellout_1_5(1);cellin_2_5(2) <= cellout_1_5(2);cellin_2_4(0) <= cellout_1_4(0);cellin_2_4(1) <= cellout_1_4(1);cellin_2_3(0) <= cellout_1_3(0);cellin_2_3(1) <= cellout_1_3(1);cellin_2_2(0) <= cellout_1_2(0);cellin_2_2(1) <= cellout_1_2(1);cellin_3_10(0) <= cellout_2_10(0);cellin_3_9(0) <= cellout_2_9(0);cellin_3_8(0) <= cellout_2_8(0);cellin_3_7(0) <= cellout_2_7(0);cellin_3_6(0) <= cellout_2_6(0);cellin_3_5(0) <= cellout_2_5(0);cellin_3_4(0) <= cellout_2_4(0);cellin_3_4(1) <= cellout_2_4(1);cellin_3_4(2) <= cellout_2_4(2);cellin_3_3(0) <= cellout_2_3(0);cellin_3_3(1) <= cellout_2_3(1);cellin_3_2(0) <= cellout_2_2(0);cellin_3_2(1) <= cellout_2_2(1);cellin_5_10(0) <= cellout_4_10(0);cellin_5_9(0) <= cellout_4_9(0);cellin_5_8(0) <= cellout_4_8(0);cellin_5_7(0) <= cellout_4_7(0);cellin_5_6(0) <= cellout_4_6(0);cellin_5_5(0) <= cellout_4_5(0);cellin_5_4(0) <= cellout_4_4(0);cellin_5_3(0) <= cellout_4_3(0);cellin_5_2(0) <= cellout_4_2(0);cellin_5_2(1) <= cellout_4_2(1);cellin_5_2(2) <= cellout_4_2(2);cellin_6_10(0) <= cellout_5_10(0);cellin_6_9(0) <= cellout_5_9(0);cellin_6_8(0) <= cellout_5_8(0);cellin_6_7(0) <= cellout_5_7(0);cellin_6_6(0) <= cellout_5_6(0);cellin_6_5(0) <= cellout_5_5(0);cellin_6_4(0) <= cellout_5_4(0);cellin_6_3(0) <= cellout_5_3(0);cellin_6_2(0) <= cellout_5_2(0);cellin_6_1(0) <= cellout_5_1(0);out_1 <= cellin_7_1;out_2 <= cellin_7_2;out_3 <= cellin_7_3;out_4 <= cellin_7_4;out_5 <= cellin_7_5;out_6 <= cellin_7_6;out_7 <= cellin_7_7;out_8 <= cellin_7_8;out_9 <= cellin_7_9;out_10 <= cellin_7_10;end generated;