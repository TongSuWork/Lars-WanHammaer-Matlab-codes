library ieee;use ieee.std_logic_1164.all;entity fir isport (  clk, reset : in std_logic;  x_0 : in std_logic_vector(5 downto 0);  y : out std_logic_vector(10 downto 0));end fir;architecture generated of fir iscomponent fir_ppport (clk, reset : in std_logic;  in_0 : in std_logic_vector(5 downto 0);  out_1_1 : out std_logic_vector(5 downto 0);  out_1_2 : out std_logic_vector(5 downto 0);  out_1_3 : out std_logic_vector(5 downto 0);  out_1_4 : out std_logic_vector(5 downto 0);  out_1_5 : out std_logic_vector(5 downto 0);  out_1_6 : out std_logic_vector(4 downto 0);  out_1_7 : out std_logic_vector(3 downto 0);  out_1_8 : out std_logic_vector(2 downto 0);  out_1_9 : out std_logic_vector(1 downto 0);  out_1_10 : out std_logic_vector(0 downto 0);  out_5_4 : out std_logic_vector(0 downto 0);  out_5_5 : out std_logic_vector(0 downto 0);  out_5_6 : out std_logic_vector(1 downto 0);  out_5_7 : out std_logic_vector(1 downto 0);  out_5_8 : out std_logic_vector(1 downto 0);  out_5_9 : out std_logic_vector(1 downto 0);  out_5_10 : out std_logic_vector(0 downto 0);  out_5_11 : out std_logic_vector(0 downto 0);  out_7_3 : out std_logic_vector(0 downto 0);  out_7_4 : out std_logic_vector(0 downto 0);  out_7_5 : out std_logic_vector(0 downto 0);  out_7_6 : out std_logic_vector(0 downto 0);  out_7_7 : out std_logic_vector(0 downto 0);  out_7_8 : out std_logic_vector(0 downto 0);  out_9_4 : out std_logic_vector(0 downto 0);  out_9_5 : out std_logic_vector(0 downto 0);  out_9_6 : out std_logic_vector(1 downto 0);  out_9_7 : out std_logic_vector(1 downto 0);  out_9_8 : out std_logic_vector(1 downto 0);  out_9_9 : out std_logic_vector(1 downto 0);  out_9_10 : out std_logic_vector(0 downto 0);  out_9_11 : out std_logic_vector(0 downto 0);  out_13_1 : out std_logic_vector(5 downto 0);  out_13_2 : out std_logic_vector(5 downto 0);  out_13_3 : out std_logic_vector(5 downto 0);  out_13_4 : out std_logic_vector(5 downto 0);  out_13_5 : out std_logic_vector(5 downto 0);  out_13_6 : out std_logic_vector(4 downto 0);  out_13_7 : out std_logic_vector(3 downto 0);  out_13_8 : out std_logic_vector(2 downto 0);  out_13_9 : out std_logic_vector(1 downto 0);  out_13_10 : out std_logic_vector(0 downto 0));end component;component fir_csport (  clk, reset : in std_logic;  in_1_1 : in std_logic_vector(5 downto 0);  in_1_2 : in std_logic_vector(5 downto 0);  in_1_3 : in std_logic_vector(5 downto 0);  in_1_4 : in std_logic_vector(5 downto 0);  in_1_5 : in std_logic_vector(5 downto 0);  in_1_6 : in std_logic_vector(4 downto 0);  in_1_7 : in std_logic_vector(3 downto 0);  in_1_8 : in std_logic_vector(2 downto 0);  in_1_9 : in std_logic_vector(1 downto 0);  in_1_10 : in std_logic_vector(0 downto 0);  in_5_4 : in std_logic_vector(0 downto 0);  in_5_5 : in std_logic_vector(0 downto 0);  in_5_6 : in std_logic_vector(1 downto 0);  in_5_7 : in std_logic_vector(1 downto 0);  in_5_8 : in std_logic_vector(1 downto 0);  in_5_9 : in std_logic_vector(1 downto 0);  in_5_10 : in std_logic_vector(0 downto 0);  in_5_11 : in std_logic_vector(0 downto 0);  in_7_3 : in std_logic_vector(0 downto 0);  in_7_4 : in std_logic_vector(0 downto 0);  in_7_5 : in std_logic_vector(0 downto 0);  in_7_6 : in std_logic_vector(0 downto 0);  in_7_7 : in std_logic_vector(0 downto 0);  in_7_8 : in std_logic_vector(0 downto 0);  in_9_4 : in std_logic_vector(0 downto 0);  in_9_5 : in std_logic_vector(0 downto 0);  in_9_6 : in std_logic_vector(1 downto 0);  in_9_7 : in std_logic_vector(1 downto 0);  in_9_8 : in std_logic_vector(1 downto 0);  in_9_9 : in std_logic_vector(1 downto 0);  in_9_10 : in std_logic_vector(0 downto 0);  in_9_11 : in std_logic_vector(0 downto 0);  in_13_1 : in std_logic_vector(5 downto 0);  in_13_2 : in std_logic_vector(5 downto 0);  in_13_3 : in std_logic_vector(5 downto 0);  in_13_4 : in std_logic_vector(5 downto 0);  in_13_5 : in std_logic_vector(5 downto 0);  in_13_6 : in std_logic_vector(4 downto 0);  in_13_7 : in std_logic_vector(3 downto 0);  in_13_8 : in std_logic_vector(2 downto 0);  in_13_9 : in std_logic_vector(1 downto 0);  in_13_10 : in std_logic_vector(0 downto 0);  out_1 : out std_logic_vector(1 downto 0);  out_2 : out std_logic_vector(1 downto 0);  out_3 : out std_logic_vector(1 downto 0);  out_4 : out std_logic_vector(1 downto 0);  out_5 : out std_logic_vector(1 downto 0);  out_6 : out std_logic_vector(1 downto 0);  out_7 : out std_logic_vector(1 downto 0);  out_8 : out std_logic_vector(0 downto 0);  out_9 : out std_logic_vector(0 downto 0);  out_10 : out std_logic_vector(0 downto 0);  out_11 : out std_logic_vector(0 downto 0));end component;component fir_vmaport (  clk, reset : in std_logic;  in_1_1 : in std_logic_vector(1 downto 0);  in_1_2 : in std_logic_vector(1 downto 0);  in_1_3 : in std_logic_vector(1 downto 0);  in_1_4 : in std_logic_vector(1 downto 0);  in_1_5 : in std_logic_vector(1 downto 0);  in_1_6 : in std_logic_vector(1 downto 0);  in_1_7 : in std_logic_vector(1 downto 0);  in_1_8 : in std_logic_vector(0 downto 0);  in_1_9 : in std_logic_vector(0 downto 0);  in_1_10 : in std_logic_vector(0 downto 0);  in_1_11 : in std_logic_vector(0 downto 0);  out_1 : out std_logic_vector(0 downto 0);  out_2 : out std_logic_vector(0 downto 0);  out_3 : out std_logic_vector(0 downto 0);  out_4 : out std_logic_vector(0 downto 0);  out_5 : out std_logic_vector(0 downto 0);  out_6 : out std_logic_vector(0 downto 0);  out_7 : out std_logic_vector(0 downto 0);  out_8 : out std_logic_vector(0 downto 0);  out_9 : out std_logic_vector(0 downto 0);  out_10 : out std_logic_vector(0 downto 0);  out_11 : out std_logic_vector(0 downto 0));end component;signal pp_1_1 : std_logic_vector(5 downto 0);signal pp_1_2 : std_logic_vector(5 downto 0);signal pp_1_3 : std_logic_vector(5 downto 0);signal pp_1_4 : std_logic_vector(5 downto 0);signal pp_1_5 : std_logic_vector(5 downto 0);signal pp_1_6 : std_logic_vector(4 downto 0);signal pp_1_7 : std_logic_vector(3 downto 0);signal pp_1_8 : std_logic_vector(2 downto 0);signal pp_1_9 : std_logic_vector(1 downto 0);signal pp_1_10 : std_logic_vector(0 downto 0);signal pp_5_4 : std_logic_vector(0 downto 0);signal pp_5_5 : std_logic_vector(0 downto 0);signal pp_5_6 : std_logic_vector(1 downto 0);signal pp_5_7 : std_logic_vector(1 downto 0);signal pp_5_8 : std_logic_vector(1 downto 0);signal pp_5_9 : std_logic_vector(1 downto 0);signal pp_5_10 : std_logic_vector(0 downto 0);signal pp_5_11 : std_logic_vector(0 downto 0);signal pp_7_3 : std_logic_vector(0 downto 0);signal pp_7_4 : std_logic_vector(0 downto 0);signal pp_7_5 : std_logic_vector(0 downto 0);signal pp_7_6 : std_logic_vector(0 downto 0);signal pp_7_7 : std_logic_vector(0 downto 0);signal pp_7_8 : std_logic_vector(0 downto 0);signal pp_9_4 : std_logic_vector(0 downto 0);signal pp_9_5 : std_logic_vector(0 downto 0);signal pp_9_6 : std_logic_vector(1 downto 0);signal pp_9_7 : std_logic_vector(1 downto 0);signal pp_9_8 : std_logic_vector(1 downto 0);signal pp_9_9 : std_logic_vector(1 downto 0);signal pp_9_10 : std_logic_vector(0 downto 0);signal pp_9_11 : std_logic_vector(0 downto 0);signal pp_13_1 : std_logic_vector(5 downto 0);signal pp_13_2 : std_logic_vector(5 downto 0);signal pp_13_3 : std_logic_vector(5 downto 0);signal pp_13_4 : std_logic_vector(5 downto 0);signal pp_13_5 : std_logic_vector(5 downto 0);signal pp_13_6 : std_logic_vector(4 downto 0);signal pp_13_7 : std_logic_vector(3 downto 0);signal pp_13_8 : std_logic_vector(2 downto 0);signal pp_13_9 : std_logic_vector(1 downto 0);signal pp_13_10 : std_logic_vector(0 downto 0);signal cs_1 : std_logic_vector(1 downto 0);signal cs_2 : std_logic_vector(1 downto 0);signal cs_3 : std_logic_vector(1 downto 0);signal cs_4 : std_logic_vector(1 downto 0);signal cs_5 : std_logic_vector(1 downto 0);signal cs_6 : std_logic_vector(1 downto 0);signal cs_7 : std_logic_vector(1 downto 0);signal cs_8 : std_logic_vector(0 downto 0);signal cs_9 : std_logic_vector(0 downto 0);signal cs_10 : std_logic_vector(0 downto 0);signal cs_11 : std_logic_vector(0 downto 0);beginpp_i: fir_pp port map(  clk => clk,  reset => reset,  in_0 => x_0,  out_1_1 => pp_1_1,  out_1_2 => pp_1_2,  out_1_3 => pp_1_3,  out_1_4 => pp_1_4,  out_1_5 => pp_1_5,  out_1_6 => pp_1_6,  out_1_7 => pp_1_7,  out_1_8 => pp_1_8,  out_1_9 => pp_1_9,  out_1_10 => pp_1_10,  out_5_4 => pp_5_4,  out_5_5 => pp_5_5,  out_5_6 => pp_5_6,  out_5_7 => pp_5_7,  out_5_8 => pp_5_8,  out_5_9 => pp_5_9,  out_5_10 => pp_5_10,  out_5_11 => pp_5_11,  out_7_3 => pp_7_3,  out_7_4 => pp_7_4,  out_7_5 => pp_7_5,  out_7_6 => pp_7_6,  out_7_7 => pp_7_7,  out_7_8 => pp_7_8,  out_9_4 => pp_9_4,  out_9_5 => pp_9_5,  out_9_6 => pp_9_6,  out_9_7 => pp_9_7,  out_9_8 => pp_9_8,  out_9_9 => pp_9_9,  out_9_10 => pp_9_10,  out_9_11 => pp_9_11,  out_13_1 => pp_13_1,  out_13_2 => pp_13_2,  out_13_3 => pp_13_3,  out_13_4 => pp_13_4,  out_13_5 => pp_13_5,  out_13_6 => pp_13_6,  out_13_7 => pp_13_7,  out_13_8 => pp_13_8,  out_13_9 => pp_13_9,  out_13_10 => pp_13_10);cs_i: fir_cs port map(  clk => clk,  reset => reset,  in_1_1 => pp_1_1,  in_1_2 => pp_1_2,  in_1_3 => pp_1_3,  in_1_4 => pp_1_4,  in_1_5 => pp_1_5,  in_1_6 => pp_1_6,  in_1_7 => pp_1_7,  in_1_8 => pp_1_8,  in_1_9 => pp_1_9,  in_1_10 => pp_1_10,  in_5_4 => pp_5_4,  in_5_5 => pp_5_5,  in_5_6 => pp_5_6,  in_5_7 => pp_5_7,  in_5_8 => pp_5_8,  in_5_9 => pp_5_9,  in_5_10 => pp_5_10,  in_5_11 => pp_5_11,  in_7_3 => pp_7_3,  in_7_4 => pp_7_4,  in_7_5 => pp_7_5,  in_7_6 => pp_7_6,  in_7_7 => pp_7_7,  in_7_8 => pp_7_8,  in_9_4 => pp_9_4,  in_9_5 => pp_9_5,  in_9_6 => pp_9_6,  in_9_7 => pp_9_7,  in_9_8 => pp_9_8,  in_9_9 => pp_9_9,  in_9_10 => pp_9_10,  in_9_11 => pp_9_11,  in_13_1 => pp_13_1,  in_13_2 => pp_13_2,  in_13_3 => pp_13_3,  in_13_4 => pp_13_4,  in_13_5 => pp_13_5,  in_13_6 => pp_13_6,  in_13_7 => pp_13_7,  in_13_8 => pp_13_8,  in_13_9 => pp_13_9,  in_13_10 => pp_13_10,  out_1 => cs_1,  out_2 => cs_2,  out_3 => cs_3,  out_4 => cs_4,  out_5 => cs_5,  out_6 => cs_6,  out_7 => cs_7,  out_8 => cs_8,  out_9 => cs_9,  out_10 => cs_10,  out_11 => cs_11);vma_i: fir_vma port map(  clk => clk,  reset => reset,  in_1_1 => cs_1,  in_1_2 => cs_2,  in_1_3 => cs_3,  in_1_4 => cs_4,  in_1_5 => cs_5,  in_1_6 => cs_6,  in_1_7 => cs_7,  in_1_8 => cs_8,  in_1_9 => cs_9,  in_1_10 => cs_10,  in_1_11 => cs_11,  out_1(0) => y(10),  out_2(0) => y(9),  out_3(0) => y(8),  out_4(0) => y(7),  out_5(0) => y(6),  out_6(0) => y(5),  out_7(0) => y(4),  out_8(0) => y(3),  out_9(0) => y(2),  out_10(0) => y(1),  out_11(0) => y(0));end generated;