library ieee;use ieee.std_logic_1164.all;entity fir_pp isport (clk, reset : in std_logic;  in_0 : in std_logic_vector(4 downto 0);  out_1_3 : out std_logic_vector(0 downto 0);  out_1_4 : out std_logic_vector(2 downto 0);  out_1_5 : out std_logic_vector(4 downto 0);  out_1_6 : out std_logic_vector(6 downto 0);  out_1_7 : out std_logic_vector(6 downto 0);  out_1_8 : out std_logic_vector(5 downto 0);  out_1_9 : out std_logic_vector(3 downto 0);  out_1_10 : out std_logic_vector(1 downto 0));end fir_pp;architecture generated of fir_pp iscomponent reggeneric (wordlength : positive);port (clk, reset : in std_logic;d : in std_logic_vector(wordlength-1 downto 0);q : out std_logic_vector(wordlength-1 downto 0));end component;signal in_0_0 : std_logic_vector(4 downto 0);signal in_0_1 : std_logic_vector(4 downto 0);signal in_0_2 : std_logic_vector(4 downto 0);signal in_0_3 : std_logic_vector(4 downto 0);signal in_0_4 : std_logic_vector(4 downto 0);signal in_0_5 : std_logic_vector(4 downto 0);signal in_0_6 : std_logic_vector(4 downto 0);beginin_0_0 <= in_0;in_d_0_1: reg generic map(5) port map(clk, reset, in_0_0, in_0_1);in_d_0_2: reg generic map(5) port map(clk, reset, in_0_1, in_0_2);in_d_0_3: reg generic map(5) port map(clk, reset, in_0_2, in_0_3);in_d_0_4: reg generic map(5) port map(clk, reset, in_0_3, in_0_4);in_d_0_5: reg generic map(5) port map(clk, reset, in_0_4, in_0_5);in_d_0_6: reg generic map(5) port map(clk, reset, in_0_5, in_0_6);out_1_3(0) <= not in_0_3(4);out_1_4(0) <= not in_0_2(4);out_1_4(1) <= in_0_3(3);out_1_4(2) <= not in_0_4(4);out_1_5(0) <= in_0_0(4);out_1_5(1) <= in_0_2(3);out_1_5(2) <= in_0_3(2);out_1_5(3) <= in_0_4(3);out_1_5(4) <= in_0_6(4);out_1_6(0) <= not in_0_0(3);out_1_6(1) <= in_0_2(2);out_1_6(2) <= not in_0_2(4);out_1_6(3) <= in_0_3(1);out_1_6(4) <= in_0_4(2);out_1_6(5) <= not in_0_4(4);out_1_6(6) <= not in_0_6(3);out_1_7(0) <= not in_0_0(2);out_1_7(1) <= in_0_2(1);out_1_7(2) <= in_0_2(3);out_1_7(3) <= in_0_3(0);out_1_7(4) <= in_0_4(1);out_1_7(5) <= in_0_4(3);out_1_7(6) <= not in_0_6(2);out_1_8(0) <= not in_0_0(1);out_1_8(1) <= in_0_2(0);out_1_8(2) <= in_0_2(2);out_1_8(3) <= in_0_4(0);out_1_8(4) <= in_0_4(2);out_1_8(5) <= not in_0_6(1);out_1_9(0) <= not in_0_0(0);out_1_9(1) <= in_0_2(1);out_1_9(2) <= in_0_4(1);out_1_9(3) <= not in_0_6(0);out_1_10(0) <= in_0_2(0);out_1_10(1) <= in_0_4(0);end generated;